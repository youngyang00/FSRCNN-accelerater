// SPDX-License-Identifier: MIT
// Copyright (c) 2025 Gwangsun Shin
module Axi4ConvCore#(
   parameter REQUANT = 172,
   parameter weight01_1_pe0 = 24'h10D3E8,
   parameter weight02_1_pe0 = 24'h7FD67F,
   parameter weight03_1_pe0 = 24'h0EB57F,
   parameter weight04_1_pe0 = 24'h807FEA,
   parameter weight05_1_pe0 = 24'h807F80,
   parameter weight06_1_pe0 = 24'h027FAB,
   parameter weight07_1_pe0 = 24'hEA487F,
   parameter weight08_1_pe0 = 24'h9519D2,
   parameter weight09_1_pe0 = 24'h027F01,
   parameter weight10_1_pe0 = 24'hCA20DC,
   parameter weight11_1_pe0 = 24'hC57F97,
   parameter weight12_1_pe0 = 24'hCD7F09,
   parameter weight13_1_pe0 = 24'h637F7F,
   parameter weight14_1_pe0 = 24'hEEBEF9,
   parameter weight15_1_pe0 = 24'h1DB5F0,
   parameter weight16_1_pe0 = 24'hCDD6D0,
   parameter weight17_1_pe0 = 24'h38E92C,
   parameter weight18_1_pe0 = 24'h68ABBF,
   parameter weight19_1_pe0 = 24'h5710CC,
   parameter weight20_1_pe0 = 24'h7F7F9A,
   parameter weight21_1_pe0 = 24'h477F7F,
   parameter weight22_1_pe0 = 24'h3E1A7F,
   parameter weight23_1_pe0 = 24'h6ACD6C,
   parameter weight24_1_pe0 = 24'h4FF380,
   parameter weight25_1_pe0 = 24'h8080DA,
   parameter weight26_1_pe0 = 24'h7F817F,
   parameter weight27_1_pe0 = 24'hCB3AE3,
   parameter weight28_1_pe0 = 24'h247F7F,
   parameter weight29_1_pe0 = 24'hF97F80,
   parameter weight30_1_pe0 = 24'h077F29,
   parameter weight31_1_pe0 = 24'h96D2A5,
   parameter weight32_1_pe0 = 24'h7FE171,
   parameter weight33_1_pe0 = 24'h7F7F19,
   parameter weight34_1_pe0 = 24'hC38030,
   parameter weight35_1_pe0 = 24'h837F12,
   parameter weight36_1_pe0 = 24'h8081C3,
   parameter weight01_2_pe0 = 24'hD97F20,
   parameter weight02_2_pe0 = 24'h318158,
   parameter weight03_2_pe0 = 24'h197F34,
   parameter weight04_2_pe0 = 24'h7FA479,
   parameter weight05_2_pe0 = 24'hA37C80,
   parameter weight06_2_pe0 = 24'h379EBB,
   parameter weight07_2_pe0 = 24'h6DCD7F,
   parameter weight08_2_pe0 = 24'h7F80DB,
   parameter weight09_2_pe0 = 24'h2D7F39,
   parameter weight10_2_pe0 = 24'hEA0380,
   parameter weight11_2_pe0 = 24'hDA7A33,
   parameter weight12_2_pe0 = 24'hEED814,
   parameter weight13_2_pe0 = 24'hEEC380,
   parameter weight14_2_pe0 = 24'hD11D25,
   parameter weight15_2_pe0 = 24'hDCE207,
   parameter weight16_2_pe0 = 24'h004D1E,
   parameter weight17_2_pe0 = 24'hC6DA06,
   parameter weight18_2_pe0 = 24'h7F28ED,
   parameter weight19_2_pe0 = 24'h7F7F7B,
   parameter weight20_2_pe0 = 24'h7F106F,
   parameter weight21_2_pe0 = 24'h7F7C7F,
   parameter weight22_2_pe0 = 24'h17C341,
   parameter weight23_2_pe0 = 24'hE825BE,
   parameter weight24_2_pe0 = 24'hF7F9C3,
   parameter weight25_2_pe0 = 24'h5E2F07,
   parameter weight26_2_pe0 = 24'h7F1027,
   parameter weight27_2_pe0 = 24'h3113E5,
   parameter weight28_2_pe0 = 24'h808080,
   parameter weight29_2_pe0 = 24'h808080,
   parameter weight30_2_pe0 = 24'h808080,
   parameter weight31_2_pe0 = 24'hA4300F,
   parameter weight32_2_pe0 = 24'hEC18F5,
   parameter weight33_2_pe0 = 24'hDFEBE2,
   parameter weight34_2_pe0 = 24'h170E1F,
   parameter weight35_2_pe0 = 24'hE51830,
   parameter weight36_2_pe0 = 24'hFE811C,
   parameter weight01_1_pe1 = 24'h2BFF2A,
   parameter weight02_1_pe1 = 24'h11CA16,
   parameter weight03_1_pe1 = 24'hEDD4EE,
   parameter weight04_1_pe1 = 24'h279FC0,
   parameter weight05_1_pe1 = 24'h001DA3,
   parameter weight06_1_pe1 = 24'h1B2B0E,
   parameter weight07_1_pe1 = 24'hCB2AED,
   parameter weight08_1_pe1 = 24'hF20BE4,
   parameter weight09_1_pe1 = 24'h2815FB,
   parameter weight10_1_pe1 = 24'h0CF6D2,
   parameter weight11_1_pe1 = 24'hD97FD8,
   parameter weight12_1_pe1 = 24'hF5E0D9,
   parameter weight13_1_pe1 = 24'h11F8F0,
   parameter weight14_1_pe1 = 24'h126D1C,
   parameter weight15_1_pe1 = 24'h1BF709,
   parameter weight16_1_pe1 = 24'h0E0A0B,
   parameter weight17_1_pe1 = 24'hD7FC05,
   parameter weight18_1_pe1 = 24'h14FA11,
   parameter weight19_1_pe1 = 24'hC4BE0A,
   parameter weight20_1_pe1 = 24'hD29211,
   parameter weight21_1_pe1 = 24'hF3072B,
   parameter weight22_1_pe1 = 24'h1FCBFD,
   parameter weight23_1_pe1 = 24'hFB7F18,
   parameter weight24_1_pe1 = 24'h1616F8,
   parameter weight25_1_pe1 = 24'hF24309,
   parameter weight26_1_pe1 = 24'hE728D3,
   parameter weight27_1_pe1 = 24'h110604,
   parameter weight28_1_pe1 = 24'h17FDDB,
   parameter weight29_1_pe1 = 24'h01F21F,
   parameter weight30_1_pe1 = 24'hF10E17,
   parameter weight31_1_pe1 = 24'hD8220D,
   parameter weight32_1_pe1 = 24'h0B2F14,
   parameter weight33_1_pe1 = 24'hF1EDF1,
   parameter weight34_1_pe1 = 24'hFC26F5,
   parameter weight35_1_pe1 = 24'hF85EFB,
   parameter weight36_1_pe1 = 24'hE6F4F0,
   parameter weight01_2_pe1 = 24'h52E6DA,
   parameter weight02_2_pe1 = 24'h572ACC,
   parameter weight03_2_pe1 = 24'h2079C8,
   parameter weight04_2_pe1 = 24'h80007F,
   parameter weight05_2_pe1 = 24'h8019BE,
   parameter weight06_2_pe1 = 24'hFCB706,
   parameter weight07_2_pe1 = 24'hE305E1,
   parameter weight08_2_pe1 = 24'hE92608,
   parameter weight09_2_pe1 = 24'hC0E903,
   parameter weight10_2_pe1 = 24'hAEE71F,
   parameter weight11_2_pe1 = 24'h2F7E1B,
   parameter weight12_2_pe1 = 24'h2DE68D,
   parameter weight13_2_pe1 = 24'h9BF3D3,
   parameter weight14_2_pe1 = 24'hC97E01,
   parameter weight15_2_pe1 = 24'hD6DEB2,
   parameter weight16_2_pe1 = 24'h2B12E8,
   parameter weight17_2_pe1 = 24'hD87FB7,
   parameter weight18_2_pe1 = 24'hFB4D7F,
   parameter weight19_2_pe1 = 24'h6EF5FA,
   parameter weight20_2_pe1 = 24'h0980E2,
   parameter weight21_2_pe1 = 24'h190DE0,
   parameter weight22_2_pe1 = 24'hE99DEC,
   parameter weight23_2_pe1 = 24'h1E0945,
   parameter weight24_2_pe1 = 24'h04E320,
   parameter weight25_2_pe1 = 24'hE742F4,
   parameter weight26_2_pe1 = 24'hCEBEC6,
   parameter weight27_2_pe1 = 24'hF6292F,
   parameter weight28_2_pe1 = 24'h00F87F,
   parameter weight29_2_pe1 = 24'h7E7F6E,
   parameter weight30_2_pe1 = 24'h1EDD80,
   parameter weight31_2_pe1 = 24'h7F561D,
   parameter weight32_2_pe1 = 24'hC7F207,
   parameter weight33_2_pe1 = 24'h1C1CFF,
   parameter weight34_2_pe1 = 24'hDD59DF,
   parameter weight35_2_pe1 = 24'h210153,
   parameter weight36_2_pe1 = 24'h21D708,
   parameter weight01_1_pe2 = 24'hC135DA,
   parameter weight02_1_pe2 = 24'h802AD2,
   parameter weight03_1_pe2 = 24'h2F41F0,
   parameter weight04_1_pe2 = 24'h7FBD4D,
   parameter weight05_1_pe2 = 24'h04E920,
   parameter weight06_1_pe2 = 24'hCCCBF6,
   parameter weight07_1_pe2 = 24'hEBF10E,
   parameter weight08_1_pe2 = 24'hDD36F2,
   parameter weight09_1_pe2 = 24'hE9EC24,
   parameter weight10_1_pe2 = 24'h0EF2F9,
   parameter weight11_1_pe2 = 24'h0A5AEF,
   parameter weight12_1_pe2 = 24'h2D0C0E,
   parameter weight13_1_pe2 = 24'h0E4CEF,
   parameter weight14_1_pe2 = 24'h134F2D,
   parameter weight15_1_pe2 = 24'hF6B91D,
   parameter weight16_1_pe2 = 24'h0607D8,
   parameter weight17_1_pe2 = 24'hBB570B,
   parameter weight18_1_pe2 = 24'hF6D7E9,
   parameter weight19_1_pe2 = 24'h2DF319,
   parameter weight20_1_pe2 = 24'hE97F12,
   parameter weight21_1_pe2 = 24'hEAD9CC,
   parameter weight22_1_pe2 = 24'h201622,
   parameter weight23_1_pe2 = 24'h0556F3,
   parameter weight24_1_pe2 = 24'hE1FDEA,
   parameter weight25_1_pe2 = 24'hFD03E8,
   parameter weight26_1_pe2 = 24'hF75B1A,
   parameter weight27_1_pe2 = 24'hF225F8,
   parameter weight28_1_pe2 = 24'h21190B,
   parameter weight29_1_pe2 = 24'hFD80A5,
   parameter weight30_1_pe2 = 24'hF71C2A,
   parameter weight31_1_pe2 = 24'hF7E1ED,
   parameter weight32_1_pe2 = 24'h1439BD,
   parameter weight33_1_pe2 = 24'h0F07F1,
   parameter weight34_1_pe2 = 24'hF4F2F6,
   parameter weight35_1_pe2 = 24'hDC540D,
   parameter weight36_1_pe2 = 24'h1BDD02,
   parameter weight01_2_pe2 = 24'hF6CB64,
   parameter weight02_2_pe2 = 24'h38F5BE,
   parameter weight03_2_pe2 = 24'hDECE24,
   parameter weight04_2_pe2 = 24'h808291,
   parameter weight05_2_pe2 = 24'hDB6228,
   parameter weight06_2_pe2 = 24'h4B06E6,
   parameter weight07_2_pe2 = 24'h2E12D2,
   parameter weight08_2_pe2 = 24'h0F5FE6,
   parameter weight09_2_pe2 = 24'h4026FF,
   parameter weight10_2_pe2 = 24'h0413FD,
   parameter weight11_2_pe2 = 24'h1A70BD,
   parameter weight12_2_pe2 = 24'hFA13E2,
   parameter weight13_2_pe2 = 24'hEC34DB,
   parameter weight14_2_pe2 = 24'h2025ED,
   parameter weight15_2_pe2 = 24'h014FF6,
   parameter weight16_2_pe2 = 24'hC7D717,
   parameter weight17_2_pe2 = 24'h0A3E27,
   parameter weight18_2_pe2 = 24'hFCE860,
   parameter weight19_2_pe2 = 24'h043CF1,
   parameter weight20_2_pe2 = 24'hF3D0ED,
   parameter weight21_2_pe2 = 24'h7FC1D3,
   parameter weight22_2_pe2 = 24'h12E4FE,
   parameter weight23_2_pe2 = 24'hFB01F9,
   parameter weight24_2_pe2 = 24'h1526AE,
   parameter weight25_2_pe2 = 24'hD125C7,
   parameter weight26_2_pe2 = 24'h45F112,
   parameter weight27_2_pe2 = 24'hE90609,
   parameter weight28_2_pe2 = 24'hF5E9D7,
   parameter weight29_2_pe2 = 24'h31270B,
   parameter weight30_2_pe2 = 24'h0C1E82,
   parameter weight31_2_pe2 = 24'hE90818,
   parameter weight32_2_pe2 = 24'hF8250D,
   parameter weight33_2_pe2 = 24'h040508,
   parameter weight34_2_pe2 = 24'h380115,
   parameter weight35_2_pe2 = 24'h3CCE52,
   parameter weight36_2_pe2 = 24'h900906,
   parameter weight01_1_pe3 = 24'h80BCFE,
   parameter weight02_1_pe3 = 24'h7F7FB3,
   parameter weight03_1_pe3 = 24'hEBC11C,
   parameter weight04_1_pe3 = 24'h547F78,
   parameter weight05_1_pe3 = 24'h808080,
   parameter weight06_1_pe3 = 24'hD47F80,
   parameter weight07_1_pe3 = 24'h2E7F1E,
   parameter weight08_1_pe3 = 24'h1A8082,
   parameter weight09_1_pe3 = 24'h807F7F,
   parameter weight10_1_pe3 = 24'h0B79E7,
   parameter weight11_1_pe3 = 24'h357FB6,
   parameter weight12_1_pe3 = 24'h5B8031,
   parameter weight13_1_pe3 = 24'hC4CB80,
   parameter weight14_1_pe3 = 24'h2B583D,
   parameter weight15_1_pe3 = 24'h11800F,
   parameter weight16_1_pe3 = 24'hF91904,
   parameter weight17_1_pe3 = 24'hF27F7F,
   parameter weight18_1_pe3 = 24'h0E807F,
   parameter weight19_1_pe3 = 24'h6E7F62,
   parameter weight20_1_pe3 = 24'hCC51EA,
   parameter weight21_1_pe3 = 24'h8F8080,
   parameter weight22_1_pe3 = 24'h1CAF7F,
   parameter weight23_1_pe3 = 24'hAC7E2A,
   parameter weight24_1_pe3 = 24'hBF040E,
   parameter weight25_1_pe3 = 24'h507EBE,
   parameter weight26_1_pe3 = 24'h54BE35,
   parameter weight27_1_pe3 = 24'hAB1CF8,
   parameter weight28_1_pe3 = 24'hFE7644,
   parameter weight29_1_pe3 = 24'h2CD59E,
   parameter weight30_1_pe3 = 24'h6D7D76,
   parameter weight31_1_pe3 = 24'h037E88,
   parameter weight32_1_pe3 = 24'hE280CB,
   parameter weight33_1_pe3 = 24'hF70B80,
   parameter weight34_1_pe3 = 24'hE780AC,
   parameter weight35_1_pe3 = 24'h807F5E,
   parameter weight36_1_pe3 = 24'h7F80B2,
   parameter weight01_2_pe3 = 24'h108041,
   parameter weight02_2_pe3 = 24'h107F21,
   parameter weight03_2_pe3 = 24'h110804,
   parameter weight04_2_pe3 = 24'hABC3A4,
   parameter weight05_2_pe3 = 24'hD3BBE9,
   parameter weight06_2_pe3 = 24'hFB1ED5,
   parameter weight07_2_pe3 = 24'hD346DC,
   parameter weight08_2_pe3 = 24'hAE7F27,
   parameter weight09_2_pe3 = 24'hADB87F,
   parameter weight10_2_pe3 = 24'hFBE60E,
   parameter weight11_2_pe3 = 24'h053FF6,
   parameter weight12_2_pe3 = 24'h17F5F0,
   parameter weight13_2_pe3 = 24'hA513DA,
   parameter weight14_2_pe3 = 24'hD324EE,
   parameter weight15_2_pe3 = 24'hCA09ED,
   parameter weight16_2_pe3 = 24'hFC1FF8,
   parameter weight17_2_pe3 = 24'h0335FB,
   parameter weight18_2_pe3 = 24'h04AF64,
   parameter weight19_2_pe3 = 24'hBEE914,
   parameter weight20_2_pe3 = 24'h120C25,
   parameter weight21_2_pe3 = 24'h019DCB,
   parameter weight22_2_pe3 = 24'hBFDBED,
   parameter weight23_2_pe3 = 24'hDF7431,
   parameter weight24_2_pe3 = 24'hD9BA56,
   parameter weight25_2_pe3 = 24'h3F09DF,
   parameter weight26_2_pe3 = 24'h4EDD25,
   parameter weight27_2_pe3 = 24'hFAFBE9,
   parameter weight28_2_pe3 = 24'hE1FE05,
   parameter weight29_2_pe3 = 24'hEB11D9,
   parameter weight30_2_pe3 = 24'h277F0D,
   parameter weight31_2_pe3 = 24'h4737D1,
   parameter weight32_2_pe3 = 24'h6526CB,
   parameter weight33_2_pe3 = 24'h1341DF,
   parameter weight34_2_pe3 = 24'h59F91F,
   parameter weight35_2_pe3 = 24'hEA0631,
   parameter weight36_2_pe3 = 24'h0CE11B,
   parameter weight01_1_pe4 = 24'hD561AD,
   parameter weight02_1_pe4 = 24'hE39151,
   parameter weight03_1_pe4 = 24'hF91136,
   parameter weight04_1_pe4 = 24'h7F7F7F,
   parameter weight05_1_pe4 = 24'h617F77,
   parameter weight06_1_pe4 = 24'hF0FC06,
   parameter weight07_1_pe4 = 24'h1DD2F0,
   parameter weight08_1_pe4 = 24'h398036,
   parameter weight09_1_pe4 = 24'h02AEE0,
   parameter weight10_1_pe4 = 24'hE1AB2B,
   parameter weight11_1_pe4 = 24'hE63122,
   parameter weight12_1_pe4 = 24'h4BFC5F,
   parameter weight13_1_pe4 = 24'h22F5FD,
   parameter weight14_1_pe4 = 24'hC97FF9,
   parameter weight15_1_pe4 = 24'hF023F0,
   parameter weight16_1_pe4 = 24'h0FE52B,
   parameter weight17_1_pe4 = 24'h1BF5DC,
   parameter weight18_1_pe4 = 24'h0AA1CB,
   parameter weight19_1_pe4 = 24'hAE150C,
   parameter weight20_1_pe4 = 24'h80F4F7,
   parameter weight21_1_pe4 = 24'hEA43FA,
   parameter weight22_1_pe4 = 24'hC4F4D4,
   parameter weight23_1_pe4 = 24'h1EF71A,
   parameter weight24_1_pe4 = 24'hFFF225,
   parameter weight25_1_pe4 = 24'h20977F,
   parameter weight26_1_pe4 = 24'h7FB8D1,
   parameter weight27_1_pe4 = 24'h2FDDE2,
   parameter weight28_1_pe4 = 24'hE72508,
   parameter weight29_1_pe4 = 24'hFD147F,
   parameter weight30_1_pe4 = 24'hF0E77F,
   parameter weight31_1_pe4 = 24'hF87603,
   parameter weight32_1_pe4 = 24'hCD4131,
   parameter weight33_1_pe4 = 24'h072F11,
   parameter weight34_1_pe4 = 24'hEB0ADA,
   parameter weight35_1_pe4 = 24'hEE34D0,
   parameter weight36_1_pe4 = 24'h081E01,
   parameter weight01_2_pe4 = 24'hE953F1,
   parameter weight02_2_pe4 = 24'h7F7FEF,
   parameter weight03_2_pe4 = 24'h5BCB23,
   parameter weight04_2_pe4 = 24'hEDA3C8,
   parameter weight05_2_pe4 = 24'hED8162,
   parameter weight06_2_pe4 = 24'hB17B04,
   parameter weight07_2_pe4 = 24'h6D7F03,
   parameter weight08_2_pe4 = 24'h7FDE03,
   parameter weight09_2_pe4 = 24'hDA7FEA,
   parameter weight10_2_pe4 = 24'hDE1032,
   parameter weight11_2_pe4 = 24'hCC7F03,
   parameter weight12_2_pe4 = 24'h837069,
   parameter weight13_2_pe4 = 24'h09ADC3,
   parameter weight14_2_pe4 = 24'hCCBB43,
   parameter weight15_2_pe4 = 24'hFE12F4,
   parameter weight16_2_pe4 = 24'h2A2BF4,
   parameter weight17_2_pe4 = 24'h37E615,
   parameter weight18_2_pe4 = 24'h255E14,
   parameter weight19_2_pe4 = 24'hF8043C,
   parameter weight20_2_pe4 = 24'h655C02,
   parameter weight21_2_pe4 = 24'h8D4BE8,
   parameter weight22_2_pe4 = 24'h31830A,
   parameter weight23_2_pe4 = 24'h257FD5,
   parameter weight24_2_pe4 = 24'hA37782,
   parameter weight25_2_pe4 = 24'hDCE9F8,
   parameter weight26_2_pe4 = 24'h748150,
   parameter weight27_2_pe4 = 24'h060EC5,
   parameter weight28_2_pe4 = 24'hEE28DD,
   parameter weight29_2_pe4 = 24'hA60B74,
   parameter weight30_2_pe4 = 24'h1B167F,
   parameter weight31_2_pe4 = 24'h167FF2,
   parameter weight32_2_pe4 = 24'h108024,
   parameter weight33_2_pe4 = 24'h1AF518,
   parameter weight34_2_pe4 = 24'h25F10C,
   parameter weight35_2_pe4 = 24'h82D9D4,
   parameter weight36_2_pe4 = 24'h17AB0F,
   parameter weight01_1_pe5 = 24'hD97F20,
   parameter weight02_1_pe5 = 24'h318158,
   parameter weight03_1_pe5 = 24'h197F34,
   parameter weight04_1_pe5 = 24'h7FA479,
   parameter weight05_1_pe5 = 24'hA37C80,
   parameter weight06_1_pe5 = 24'h379EBB,
   parameter weight07_1_pe5 = 24'h6DCD7F,
   parameter weight08_1_pe5 = 24'h7F80DB,
   parameter weight09_1_pe5 = 24'h2D7F39,
   parameter weight10_1_pe5 = 24'hEA0380,
   parameter weight11_1_pe5 = 24'hDA7A33,
   parameter weight12_1_pe5 = 24'hEED814,
   parameter weight13_1_pe5 = 24'hEEC380,
   parameter weight14_1_pe5 = 24'hD11D25,
   parameter weight15_1_pe5 = 24'hDCE207,
   parameter weight16_1_pe5 = 24'h004D1E,
   parameter weight17_1_pe5 = 24'hC6DA06,
   parameter weight18_1_pe5 = 24'h7F28ED,
   parameter weight19_1_pe5 = 24'h7F7F7B,
   parameter weight20_1_pe5 = 24'h7F106F,
   parameter weight21_1_pe5 = 24'h7F7C7F,
   parameter weight22_1_pe5 = 24'h17C341,
   parameter weight23_1_pe5 = 24'hE825BE,
   parameter weight24_1_pe5 = 24'hF7F9C3,
   parameter weight25_1_pe5 = 24'h5E2F07,
   parameter weight26_1_pe5 = 24'h7F1027,
   parameter weight27_1_pe5 = 24'h3113E5,
   parameter weight28_1_pe5 = 24'h808080,
   parameter weight29_1_pe5 = 24'h808080,
   parameter weight30_1_pe5 = 24'h808080,
   parameter weight31_1_pe5 = 24'hA4300F,
   parameter weight32_1_pe5 = 24'hEC18F5,
   parameter weight33_1_pe5 = 24'hDFEBE2,
   parameter weight34_1_pe5 = 24'h170E1F,
   parameter weight35_1_pe5 = 24'hE51830,
   parameter weight36_1_pe5 = 24'hFE811C,
   parameter weight01_2_pe5 = 24'h2616DA,
   parameter weight02_2_pe5 = 24'h7F800D,
   parameter weight03_2_pe5 = 24'h64EBF2,
   parameter weight04_2_pe5 = 24'h29F0F9,
   parameter weight05_2_pe5 = 24'h7F78EF,
   parameter weight06_2_pe5 = 24'h80FEF4,
   parameter weight07_2_pe5 = 24'hFDBFF9,
   parameter weight08_2_pe5 = 24'h7F070E,
   parameter weight09_2_pe5 = 24'h9F0300,
   parameter weight10_2_pe5 = 24'hEAB920,
   parameter weight11_2_pe5 = 24'h817F80,
   parameter weight12_2_pe5 = 24'h80370F,
   parameter weight13_2_pe5 = 24'hBB7FA5,
   parameter weight14_2_pe5 = 24'h80D363,
   parameter weight15_2_pe5 = 24'h80FA80,
   parameter weight16_2_pe5 = 24'h0AFCDB,
   parameter weight17_2_pe5 = 24'hAC7F1F,
   parameter weight18_2_pe5 = 24'h808009,
   parameter weight19_2_pe5 = 24'h98FBF4,
   parameter weight20_2_pe5 = 24'h8080FB,
   parameter weight21_2_pe5 = 24'h7F80EF,
   parameter weight22_2_pe5 = 24'h7FD21D,
   parameter weight23_2_pe5 = 24'h1D285D,
   parameter weight24_2_pe5 = 24'h8262C3,
   parameter weight25_2_pe5 = 24'h801403,
   parameter weight26_2_pe5 = 24'h80C60A,
   parameter weight27_2_pe5 = 24'h807FCC,
   parameter weight28_2_pe5 = 24'h2C080E,
   parameter weight29_2_pe5 = 24'h437FE1,
   parameter weight30_2_pe5 = 24'h8080F5,
   parameter weight31_2_pe5 = 24'hC46BE3,
   parameter weight32_2_pe5 = 24'h823AFB,
   parameter weight33_2_pe5 = 24'h7BE751,
   parameter weight34_2_pe5 = 24'hDB361C,
   parameter weight35_2_pe5 = 24'h7F7F35,
   parameter weight36_2_pe5 = 24'h7F9200
   
)(
   input          i_clk,
   input          i_rstn,
   output         s_axis_tready,
   input          s_axis_tvalid,
   input  [95:0]  s_axis_tdata, /* MSB: Ch12 ~ LSB:CH0 */
   output [95:0]  m_axis_tdata,
   output         m_axis_tvalid,
   input          m_axis_tready,
   output         EOL,
   output         EOF
);
localparam PE_DELAY = 11;
wire                    clr;
wire [2:0]              addr;
wire  [287:0]           Distributor_data_packed;   
wire  [7:0]             PE_Array [0:5];
wire                    Distributor_out_valid;
reg   [PE_DELAY-1:0]    Distributor_out_valid_inter;
wire  [5:0]             PE_valid_out;
wire                    PE_total_valid = &PE_valid_out & Distributor_out_valid_inter[8];
reg   [95:0]            Packed_outPixel;
reg   subCnt;
reg   backBuffer_inValid;
wire  backBuffer_prog_full;
wire  backBuffer_s_ready;
integer i;

always @(posedge i_clk) begin
   if (!i_rstn) begin
      subCnt <= 'd0;
   end
   else begin
      backBuffer_inValid <= PE_total_valid & subCnt;
      if (PE_total_valid) begin
         Packed_outPixel[95:48] <= {PE_Array[5],PE_Array[4],PE_Array[3],PE_Array[2],PE_Array[1],PE_Array[0]};
         Packed_outPixel[47:0] <= Packed_outPixel[95:48];
         subCnt <= subCnt + 'd1;
      end
   end
end

always @(posedge i_clk) begin
   Distributor_out_valid_inter[0] <= Distributor_out_valid;
   for (i = 0; i < PE_DELAY - 1; i = i + 1) begin
      Distributor_out_valid_inter[i + 1] <= Distributor_out_valid_inter[i];
   end
end

AxiBramDistributor Distributor(
   .i_clk(i_clk), //input             
   .i_rstn(i_rstn), //input             
   .s_axis_tready(s_axis_tready), //output         
   .s_axis_tvalid(s_axis_tvalid), //input             
   .s_axis_tdata(s_axis_tdata), //input [95:0]      
   .i_backBuffer_prog_full(backBuffer_prog_full),
   .i_backBuffer_s_ready(backBuffer_s_ready),
   .o_data_packed(Distributor_data_packed), //output   [287:0]  
   .o_clr(clr), //output            
   .o_addr(addr), //output [2:0]   
   .o_valid(Distributor_out_valid)
);

fifo_generator_0 backBuffer(
  .s_aclk(i_clk),                  // input wire s_aclk
  .s_aresetn(i_rstn),            // input wire s_aresetn
  .s_axis_tvalid(backBuffer_inValid),    // input wire s_axis_tvalid
  .s_axis_tready(backBuffer_s_ready),    // output wire s_axis_tready
  .s_axis_tdata({{32'b0},Packed_outPixel}),      // input wire [127 : 0] s_axis_tdata
  .s_axis_tuser(),      // input wire [3 : 0] s_axis_tuser
  .m_axis_tvalid(m_axis_tvalid),    // output wire m_axis_tvalid
  .m_axis_tready(m_axis_tready),    // input wire m_axis_tready
  .m_axis_tdata(m_axis_tdata),      // output wire [127 : 0] m_axis_tdata
  .m_axis_tuser(),      // output wire [3 : 0] m_axis_tuser
  .axis_prog_full(backBuffer_prog_full)  // output wire axis_prog_full
);

PE_Array#(
   .REQUANT(REQUANT),
   .weight01_1(weight01_1_pe0),
   .weight02_1(weight02_1_pe0),
   .weight03_1(weight03_1_pe0),
   .weight04_1(weight04_1_pe0),
   .weight05_1(weight05_1_pe0),
   .weight06_1(weight06_1_pe0),
   .weight07_1(weight07_1_pe0),
   .weight08_1(weight08_1_pe0),
   .weight09_1(weight09_1_pe0),
   .weight10_1(weight10_1_pe0),
   .weight11_1(weight11_1_pe0),
   .weight12_1(weight12_1_pe0),
   .weight13_1(weight13_1_pe0),
   .weight14_1(weight14_1_pe0),
   .weight15_1(weight15_1_pe0),
   .weight16_1(weight16_1_pe0),
   .weight17_1(weight17_1_pe0),
   .weight18_1(weight18_1_pe0),
   .weight19_1(weight19_1_pe0),
   .weight20_1(weight20_1_pe0),
   .weight21_1(weight21_1_pe0),
   .weight22_1(weight22_1_pe0),
   .weight23_1(weight23_1_pe0),
   .weight24_1(weight24_1_pe0),
   .weight25_1(weight25_1_pe0),
   .weight26_1(weight26_1_pe0),
   .weight27_1(weight27_1_pe0),
   .weight28_1(weight28_1_pe0),
   .weight29_1(weight29_1_pe0),
   .weight30_1(weight30_1_pe0),
   .weight31_1(weight31_1_pe0),
   .weight32_1(weight32_1_pe0),
   .weight33_1(weight33_1_pe0),
   .weight34_1(weight34_1_pe0),
   .weight35_1(weight35_1_pe0),
   .weight36_1(weight36_1_pe0),
   .weight01_2(weight01_2_pe0),
   .weight02_2(weight02_2_pe0),
   .weight03_2(weight03_2_pe0),
   .weight04_2(weight04_2_pe0),
   .weight05_2(weight05_2_pe0),
   .weight06_2(weight06_2_pe0),
   .weight07_2(weight07_2_pe0),
   .weight08_2(weight08_2_pe0),
   .weight09_2(weight09_2_pe0),
   .weight10_2(weight10_2_pe0),
   .weight11_2(weight11_2_pe0),
   .weight12_2(weight12_2_pe0),
   .weight13_2(weight13_2_pe0),
   .weight14_2(weight14_2_pe0),
   .weight15_2(weight15_2_pe0),
   .weight16_2(weight16_2_pe0),
   .weight17_2(weight17_2_pe0),
   .weight18_2(weight18_2_pe0),
   .weight19_2(weight19_2_pe0),
   .weight20_2(weight20_2_pe0),
   .weight21_2(weight21_2_pe0),
   .weight22_2(weight22_2_pe0),
   .weight23_2(weight23_2_pe0),
   .weight24_2(weight24_2_pe0),
   .weight25_2(weight25_2_pe0),
   .weight26_2(weight26_2_pe0),
   .weight27_2(weight27_2_pe0),
   .weight28_2(weight28_2_pe0),
   .weight29_2(weight29_2_pe0),
   .weight30_2(weight30_2_pe0),
   .weight31_2(weight31_2_pe0),
   .weight32_2(weight32_2_pe0),
   .weight33_2(weight33_2_pe0),
   .weight34_2(weight34_2_pe0),
   .weight35_2(weight35_2_pe0),
   .weight36_2(weight36_2_pe0)
)pe_array0(
   .i_clk(i_clk), //input                
   .i_clr(clr), //input                
   .i_en(1'b1), //input                
   .i_addr(addr), //input       [2:0]    
   .i_pixel(Distributor_data_packed),  //input       [287:0]  
   .o_valid(PE_valid_out[0]), //output            
   .o_result(PE_Array[0]) //output   [7:0]    
);

PE_Array#(
   .REQUANT(REQUANT),
   .weight01_1(weight01_1_pe1),
   .weight02_1(weight02_1_pe1),
   .weight03_1(weight03_1_pe1),
   .weight04_1(weight04_1_pe1),
   .weight05_1(weight05_1_pe1),
   .weight06_1(weight06_1_pe1),
   .weight07_1(weight07_1_pe1),
   .weight08_1(weight08_1_pe1),
   .weight09_1(weight09_1_pe1),
   .weight10_1(weight10_1_pe1),
   .weight11_1(weight11_1_pe1),
   .weight12_1(weight12_1_pe1),
   .weight13_1(weight13_1_pe1),
   .weight14_1(weight14_1_pe1),
   .weight15_1(weight15_1_pe1),
   .weight16_1(weight16_1_pe1),
   .weight17_1(weight17_1_pe1),
   .weight18_1(weight18_1_pe1),
   .weight19_1(weight19_1_pe1),
   .weight20_1(weight20_1_pe1),
   .weight21_1(weight21_1_pe1),
   .weight22_1(weight22_1_pe1),
   .weight23_1(weight23_1_pe1),
   .weight24_1(weight24_1_pe1),
   .weight25_1(weight25_1_pe1),
   .weight26_1(weight26_1_pe1),
   .weight27_1(weight27_1_pe1),
   .weight28_1(weight28_1_pe1),
   .weight29_1(weight29_1_pe1),
   .weight30_1(weight30_1_pe1),
   .weight31_1(weight31_1_pe1),
   .weight32_1(weight32_1_pe1),
   .weight33_1(weight33_1_pe1),
   .weight34_1(weight34_1_pe1),
   .weight35_1(weight35_1_pe1),
   .weight36_1(weight36_1_pe1),
   .weight01_2(weight01_2_pe1),
   .weight02_2(weight02_2_pe1),
   .weight03_2(weight03_2_pe1),
   .weight04_2(weight04_2_pe1),
   .weight05_2(weight05_2_pe1),
   .weight06_2(weight06_2_pe1),
   .weight07_2(weight07_2_pe1),
   .weight08_2(weight08_2_pe1),
   .weight09_2(weight09_2_pe1),
   .weight10_2(weight10_2_pe1),
   .weight11_2(weight11_2_pe1),
   .weight12_2(weight12_2_pe1),
   .weight13_2(weight13_2_pe1),
   .weight14_2(weight14_2_pe1),
   .weight15_2(weight15_2_pe1),
   .weight16_2(weight16_2_pe1),
   .weight17_2(weight17_2_pe1),
   .weight18_2(weight18_2_pe1),
   .weight19_2(weight19_2_pe1),
   .weight20_2(weight20_2_pe1),
   .weight21_2(weight21_2_pe1),
   .weight22_2(weight22_2_pe1),
   .weight23_2(weight23_2_pe1),
   .weight24_2(weight24_2_pe1),
   .weight25_2(weight25_2_pe1),
   .weight26_2(weight26_2_pe1),
   .weight27_2(weight27_2_pe1),
   .weight28_2(weight28_2_pe1),
   .weight29_2(weight29_2_pe1),
   .weight30_2(weight30_2_pe1),
   .weight31_2(weight31_2_pe1),
   .weight32_2(weight32_2_pe1),
   .weight33_2(weight33_2_pe1),
   .weight34_2(weight34_2_pe1),
   .weight35_2(weight35_2_pe1),
   .weight36_2(weight36_2_pe1)
)pe_array1(
   .i_clk(i_clk), //input                
   .i_clr(clr), //input                
   .i_en(1'b1), //input                
   .i_addr(addr), //input       [2:0]    
   .i_pixel(Distributor_data_packed),  //input       [287:0]  
   .o_valid(PE_valid_out[1]), //output            
   .o_result(PE_Array[1]) //output   [7:0]    
);

PE_Array#(
   .REQUANT(REQUANT),
   .weight01_1(weight01_1_pe2),
   .weight02_1(weight02_1_pe2),
   .weight03_1(weight03_1_pe2),
   .weight04_1(weight04_1_pe2),
   .weight05_1(weight05_1_pe2),
   .weight06_1(weight06_1_pe2),
   .weight07_1(weight07_1_pe2),
   .weight08_1(weight08_1_pe2),
   .weight09_1(weight09_1_pe2),
   .weight10_1(weight10_1_pe2),
   .weight11_1(weight11_1_pe2),
   .weight12_1(weight12_1_pe2),
   .weight13_1(weight13_1_pe2),
   .weight14_1(weight14_1_pe2),
   .weight15_1(weight15_1_pe2),
   .weight16_1(weight16_1_pe2),
   .weight17_1(weight17_1_pe2),
   .weight18_1(weight18_1_pe2),
   .weight19_1(weight19_1_pe2),
   .weight20_1(weight20_1_pe2),
   .weight21_1(weight21_1_pe2),
   .weight22_1(weight22_1_pe2),
   .weight23_1(weight23_1_pe2),
   .weight24_1(weight24_1_pe2),
   .weight25_1(weight25_1_pe2),
   .weight26_1(weight26_1_pe2),
   .weight27_1(weight27_1_pe2),
   .weight28_1(weight28_1_pe2),
   .weight29_1(weight29_1_pe2),
   .weight30_1(weight30_1_pe2),
   .weight31_1(weight31_1_pe2),
   .weight32_1(weight32_1_pe2),
   .weight33_1(weight33_1_pe2),
   .weight34_1(weight34_1_pe2),
   .weight35_1(weight35_1_pe2),
   .weight36_1(weight36_1_pe2),
   .weight01_2(weight01_2_pe2),
   .weight02_2(weight02_2_pe2),
   .weight03_2(weight03_2_pe2),
   .weight04_2(weight04_2_pe2),
   .weight05_2(weight05_2_pe2),
   .weight06_2(weight06_2_pe2),
   .weight07_2(weight07_2_pe2),
   .weight08_2(weight08_2_pe2),
   .weight09_2(weight09_2_pe2),
   .weight10_2(weight10_2_pe2),
   .weight11_2(weight11_2_pe2),
   .weight12_2(weight12_2_pe2),
   .weight13_2(weight13_2_pe2),
   .weight14_2(weight14_2_pe2),
   .weight15_2(weight15_2_pe2),
   .weight16_2(weight16_2_pe2),
   .weight17_2(weight17_2_pe2),
   .weight18_2(weight18_2_pe2),
   .weight19_2(weight19_2_pe2),
   .weight20_2(weight20_2_pe2),
   .weight21_2(weight21_2_pe2),
   .weight22_2(weight22_2_pe2),
   .weight23_2(weight23_2_pe2),
   .weight24_2(weight24_2_pe2),
   .weight25_2(weight25_2_pe2),
   .weight26_2(weight26_2_pe2),
   .weight27_2(weight27_2_pe2),
   .weight28_2(weight28_2_pe2),
   .weight29_2(weight29_2_pe2),
   .weight30_2(weight30_2_pe2),
   .weight31_2(weight31_2_pe2),
   .weight32_2(weight32_2_pe2),
   .weight33_2(weight33_2_pe2),
   .weight34_2(weight34_2_pe2),
   .weight35_2(weight35_2_pe2),
   .weight36_2(weight36_2_pe2)
)pe_array2(
   .i_clk(i_clk), //input                
   .i_clr(clr), //input                
   .i_en(1'b1), //input                
   .i_addr(addr), //input       [2:0]    
   .i_pixel(Distributor_data_packed),  //input       [287:0]  
   .o_valid(PE_valid_out[2]), //output            
   .o_result(PE_Array[2]) //output   [7:0]    
);

PE_Array#(
   .REQUANT(REQUANT),
   .weight01_1(weight01_1_pe3),
   .weight02_1(weight02_1_pe3),
   .weight03_1(weight03_1_pe3),
   .weight04_1(weight04_1_pe3),
   .weight05_1(weight05_1_pe3),
   .weight06_1(weight06_1_pe3),
   .weight07_1(weight07_1_pe3),
   .weight08_1(weight08_1_pe3),
   .weight09_1(weight09_1_pe3),
   .weight10_1(weight10_1_pe3),
   .weight11_1(weight11_1_pe3),
   .weight12_1(weight12_1_pe3),
   .weight13_1(weight13_1_pe3),
   .weight14_1(weight14_1_pe3),
   .weight15_1(weight15_1_pe3),
   .weight16_1(weight16_1_pe3),
   .weight17_1(weight17_1_pe3),
   .weight18_1(weight18_1_pe3),
   .weight19_1(weight19_1_pe3),
   .weight20_1(weight20_1_pe3),
   .weight21_1(weight21_1_pe3),
   .weight22_1(weight22_1_pe3),
   .weight23_1(weight23_1_pe3),
   .weight24_1(weight24_1_pe3),
   .weight25_1(weight25_1_pe3),
   .weight26_1(weight26_1_pe3),
   .weight27_1(weight27_1_pe3),
   .weight28_1(weight28_1_pe3),
   .weight29_1(weight29_1_pe3),
   .weight30_1(weight30_1_pe3),
   .weight31_1(weight31_1_pe3),
   .weight32_1(weight32_1_pe3),
   .weight33_1(weight33_1_pe3),
   .weight34_1(weight34_1_pe3),
   .weight35_1(weight35_1_pe3),
   .weight36_1(weight36_1_pe3),
   .weight01_2(weight01_2_pe3),
   .weight02_2(weight02_2_pe3),
   .weight03_2(weight03_2_pe3),
   .weight04_2(weight04_2_pe3),
   .weight05_2(weight05_2_pe3),
   .weight06_2(weight06_2_pe3),
   .weight07_2(weight07_2_pe3),
   .weight08_2(weight08_2_pe3),
   .weight09_2(weight09_2_pe3),
   .weight10_2(weight10_2_pe3),
   .weight11_2(weight11_2_pe3),
   .weight12_2(weight12_2_pe3),
   .weight13_2(weight13_2_pe3),
   .weight14_2(weight14_2_pe3),
   .weight15_2(weight15_2_pe3),
   .weight16_2(weight16_2_pe3),
   .weight17_2(weight17_2_pe3),
   .weight18_2(weight18_2_pe3),
   .weight19_2(weight19_2_pe3),
   .weight20_2(weight20_2_pe3),
   .weight21_2(weight21_2_pe3),
   .weight22_2(weight22_2_pe3),
   .weight23_2(weight23_2_pe3),
   .weight24_2(weight24_2_pe3),
   .weight25_2(weight25_2_pe3),
   .weight26_2(weight26_2_pe3),
   .weight27_2(weight27_2_pe3),
   .weight28_2(weight28_2_pe3),
   .weight29_2(weight29_2_pe3),
   .weight30_2(weight30_2_pe3),
   .weight31_2(weight31_2_pe3),
   .weight32_2(weight32_2_pe3),
   .weight33_2(weight33_2_pe3),
   .weight34_2(weight34_2_pe3),
   .weight35_2(weight35_2_pe3),
   .weight36_2(weight36_2_pe3)
)pe_array3(
   .i_clk(i_clk), //input                
   .i_clr(clr), //input                
   .i_en(1'b1), //input                
   .i_addr(addr), //input       [2:0]    
   .i_pixel(Distributor_data_packed),  //input       [287:0]  
   .o_valid(PE_valid_out[3]), //output            
   .o_result(PE_Array[3]) //output   [7:0]    
);

PE_Array#(
   .REQUANT(REQUANT),
   .weight01_1(weight01_1_pe4),
   .weight02_1(weight02_1_pe4),
   .weight03_1(weight03_1_pe4),
   .weight04_1(weight04_1_pe4),
   .weight05_1(weight05_1_pe4),
   .weight06_1(weight06_1_pe4),
   .weight07_1(weight07_1_pe4),
   .weight08_1(weight08_1_pe4),
   .weight09_1(weight09_1_pe4),
   .weight10_1(weight10_1_pe4),
   .weight11_1(weight11_1_pe4),
   .weight12_1(weight12_1_pe4),
   .weight13_1(weight13_1_pe4),
   .weight14_1(weight14_1_pe4),
   .weight15_1(weight15_1_pe4),
   .weight16_1(weight16_1_pe4),
   .weight17_1(weight17_1_pe4),
   .weight18_1(weight18_1_pe4),
   .weight19_1(weight19_1_pe4),
   .weight20_1(weight20_1_pe4),
   .weight21_1(weight21_1_pe4),
   .weight22_1(weight22_1_pe4),
   .weight23_1(weight23_1_pe4),
   .weight24_1(weight24_1_pe4),
   .weight25_1(weight25_1_pe4),
   .weight26_1(weight26_1_pe4),
   .weight27_1(weight27_1_pe4),
   .weight28_1(weight28_1_pe4),
   .weight29_1(weight29_1_pe4),
   .weight30_1(weight30_1_pe4),
   .weight31_1(weight31_1_pe4),
   .weight32_1(weight32_1_pe4),
   .weight33_1(weight33_1_pe4),
   .weight34_1(weight34_1_pe4),
   .weight35_1(weight35_1_pe4),
   .weight36_1(weight36_1_pe4),
   .weight01_2(weight01_2_pe4),
   .weight02_2(weight02_2_pe4),
   .weight03_2(weight03_2_pe4),
   .weight04_2(weight04_2_pe4),
   .weight05_2(weight05_2_pe4),
   .weight06_2(weight06_2_pe4),
   .weight07_2(weight07_2_pe4),
   .weight08_2(weight08_2_pe4),
   .weight09_2(weight09_2_pe4),
   .weight10_2(weight10_2_pe4),
   .weight11_2(weight11_2_pe4),
   .weight12_2(weight12_2_pe4),
   .weight13_2(weight13_2_pe4),
   .weight14_2(weight14_2_pe4),
   .weight15_2(weight15_2_pe4),
   .weight16_2(weight16_2_pe4),
   .weight17_2(weight17_2_pe4),
   .weight18_2(weight18_2_pe4),
   .weight19_2(weight19_2_pe4),
   .weight20_2(weight20_2_pe4),
   .weight21_2(weight21_2_pe4),
   .weight22_2(weight22_2_pe4),
   .weight23_2(weight23_2_pe4),
   .weight24_2(weight24_2_pe4),
   .weight25_2(weight25_2_pe4),
   .weight26_2(weight26_2_pe4),
   .weight27_2(weight27_2_pe4),
   .weight28_2(weight28_2_pe4),
   .weight29_2(weight29_2_pe4),
   .weight30_2(weight30_2_pe4),
   .weight31_2(weight31_2_pe4),
   .weight32_2(weight32_2_pe4),
   .weight33_2(weight33_2_pe4),
   .weight34_2(weight34_2_pe4),
   .weight35_2(weight35_2_pe4),
   .weight36_2(weight36_2_pe4)
)pe_array4(
   .i_clk(i_clk), //input                
   .i_clr(clr), //input                
   .i_en(1'b1), //input                
   .i_addr(addr), //input       [2:0]    
   .i_pixel(Distributor_data_packed),  //input       [287:0]  
   .o_valid(PE_valid_out[4]), //output            
   .o_result(PE_Array[4]) //output   [7:0]    
);

PE_Array#(
   .REQUANT(REQUANT),
   .weight01_1(weight01_1_pe5),
   .weight02_1(weight02_1_pe5),
   .weight03_1(weight03_1_pe5),
   .weight04_1(weight04_1_pe5),
   .weight05_1(weight05_1_pe5),
   .weight06_1(weight06_1_pe5),
   .weight07_1(weight07_1_pe5),
   .weight08_1(weight08_1_pe5),
   .weight09_1(weight09_1_pe5),
   .weight10_1(weight10_1_pe5),
   .weight11_1(weight11_1_pe5),
   .weight12_1(weight12_1_pe5),
   .weight13_1(weight13_1_pe5),
   .weight14_1(weight14_1_pe5),
   .weight15_1(weight15_1_pe5),
   .weight16_1(weight16_1_pe5),
   .weight17_1(weight17_1_pe5),
   .weight18_1(weight18_1_pe5),
   .weight19_1(weight19_1_pe5),
   .weight20_1(weight20_1_pe5),
   .weight21_1(weight21_1_pe5),
   .weight22_1(weight22_1_pe5),
   .weight23_1(weight23_1_pe5),
   .weight24_1(weight24_1_pe5),
   .weight25_1(weight25_1_pe5),
   .weight26_1(weight26_1_pe5),
   .weight27_1(weight27_1_pe5),
   .weight28_1(weight28_1_pe5),
   .weight29_1(weight29_1_pe5),
   .weight30_1(weight30_1_pe5),
   .weight31_1(weight31_1_pe5),
   .weight32_1(weight32_1_pe5),
   .weight33_1(weight33_1_pe5),
   .weight34_1(weight34_1_pe5),
   .weight35_1(weight35_1_pe5),
   .weight36_1(weight36_1_pe5),
   .weight01_2(weight01_2_pe5),
   .weight02_2(weight02_2_pe5),
   .weight03_2(weight03_2_pe5),
   .weight04_2(weight04_2_pe5),
   .weight05_2(weight05_2_pe5),
   .weight06_2(weight06_2_pe5),
   .weight07_2(weight07_2_pe5),
   .weight08_2(weight08_2_pe5),
   .weight09_2(weight09_2_pe5),
   .weight10_2(weight10_2_pe5),
   .weight11_2(weight11_2_pe5),
   .weight12_2(weight12_2_pe5),
   .weight13_2(weight13_2_pe5),
   .weight14_2(weight14_2_pe5),
   .weight15_2(weight15_2_pe5),
   .weight16_2(weight16_2_pe5),
   .weight17_2(weight17_2_pe5),
   .weight18_2(weight18_2_pe5),
   .weight19_2(weight19_2_pe5),
   .weight20_2(weight20_2_pe5),
   .weight21_2(weight21_2_pe5),
   .weight22_2(weight22_2_pe5),
   .weight23_2(weight23_2_pe5),
   .weight24_2(weight24_2_pe5),
   .weight25_2(weight25_2_pe5),
   .weight26_2(weight26_2_pe5),
   .weight27_2(weight27_2_pe5),
   .weight28_2(weight28_2_pe5),
   .weight29_2(weight29_2_pe5),
   .weight30_2(weight30_2_pe5),
   .weight31_2(weight31_2_pe5),
   .weight32_2(weight32_2_pe5),
   .weight33_2(weight33_2_pe5),
   .weight34_2(weight34_2_pe5),
   .weight35_2(weight35_2_pe5),
   .weight36_2(weight36_2_pe5)
)pe_array5(
   .i_clk(i_clk), //input                
   .i_clr(clr), //input                
   .i_en(1'b1), //input                
   .i_addr(addr), //input       [2:0]    
   .i_pixel(Distributor_data_packed),  //input       [287:0]  
   .o_valid(PE_valid_out[5]), //output            
   .o_result(PE_Array[5]) //output   [7:0]    
);

endmodule