module AxiMappingLayer(
   input          i_clk,
   input          i_rstn,
   input  [95:0]  s_axis_tdata,
   input          s_axis_tvalid,
   output         s_axis_tready,
   output [95:0]  m_axis_tdata,
   output         m_axis_tvalid,
   input          m_axis_tready,
   output         EOL,
   output         EOF
);

reg [8:0] outXcnt;
reg [7:0] outYcnt;

assign EOL = (outXcnt == 'd319) & m_axis_tvalid;
assign EOF = ((outXcnt == 'd319) & (outYcnt == 'd179)) & m_axis_tvalid;
always @(posedge i_clk) begin
   if (!i_rstn) begin
      outXcnt <= 'd0;
      outYcnt <= 'd0;
   end
   else begin
      if (m_axis_tvalid & m_axis_tready) begin
         if (outXcnt == 'd319) begin
            outXcnt <= 'd0;
            if(outYcnt == 'd179)begin
               outYcnt <= 'd0;
            end
            else begin 
               outYcnt <= outYcnt + 'd1;
            end
         end
         else begin
            outXcnt <= outXcnt + 'd1;
         end
      end
   end
end

wire [95:0] m_axis_tdata_core [0:2];
wire        m_axis_tvalid_core [0:2];
wire        m_axis_tready_core [0:2];

Axi4ConvCore#(
   .REQUANT(172),
   .weight01_1_pe0(24'h10D3E8),
   .weight02_1_pe0(24'h7FD67F),
   .weight03_1_pe0(24'h0EB57F),
   .weight04_1_pe0(24'h807FEA),
   .weight05_1_pe0(24'h807F80),
   .weight06_1_pe0(24'h027FAB),
   .weight07_1_pe0(24'hEA487F),
   .weight08_1_pe0(24'h9519D2),
   .weight09_1_pe0(24'h027F01),
   .weight10_1_pe0(24'hCA20DC),
   .weight11_1_pe0(24'hC57F97),
   .weight12_1_pe0(24'hCD7F09),
   .weight13_1_pe0(24'h637F7F),
   .weight14_1_pe0(24'hEEBEF9),
   .weight15_1_pe0(24'h1DB5F0),
   .weight16_1_pe0(24'hCDD6D0),
   .weight17_1_pe0(24'h38E92C),
   .weight18_1_pe0(24'h68ABBF),
   .weight19_1_pe0(24'h5710CC),
   .weight20_1_pe0(24'h7F7F9A),
   .weight21_1_pe0(24'h477F7F),
   .weight22_1_pe0(24'h3E1A7F),
   .weight23_1_pe0(24'h6ACD6C),
   .weight24_1_pe0(24'h4FF380),
   .weight25_1_pe0(24'h8080DA),
   .weight26_1_pe0(24'h7F817F),
   .weight27_1_pe0(24'hCB3AE3),
   .weight28_1_pe0(24'h247F7F),
   .weight29_1_pe0(24'hF97F80),
   .weight30_1_pe0(24'h077F29),
   .weight31_1_pe0(24'h96D2A5),
   .weight32_1_pe0(24'h7FE171),
   .weight33_1_pe0(24'h7F7F19),
   .weight34_1_pe0(24'hC38030),
   .weight35_1_pe0(24'h837F12),
   .weight36_1_pe0(24'h8081C3),
   .weight01_2_pe0(24'hD97F20),
   .weight02_2_pe0(24'h318158),
   .weight03_2_pe0(24'h197F34),
   .weight04_2_pe0(24'h7FA479),
   .weight05_2_pe0(24'hA37C80),
   .weight06_2_pe0(24'h379EBB),
   .weight07_2_pe0(24'h6DCD7F),
   .weight08_2_pe0(24'h7F80DB),
   .weight09_2_pe0(24'h2D7F39),
   .weight10_2_pe0(24'hEA0380),
   .weight11_2_pe0(24'hDA7A33),
   .weight12_2_pe0(24'hEED814),
   .weight13_2_pe0(24'hEEC380),
   .weight14_2_pe0(24'hD11D25),
   .weight15_2_pe0(24'hDCE207),
   .weight16_2_pe0(24'h004D1E),
   .weight17_2_pe0(24'hC6DA06),
   .weight18_2_pe0(24'h7F28ED),
   .weight19_2_pe0(24'h7F7F7B),
   .weight20_2_pe0(24'h7F106F),
   .weight21_2_pe0(24'h7F7C7F),
   .weight22_2_pe0(24'h17C341),
   .weight23_2_pe0(24'hE825BE),
   .weight24_2_pe0(24'hF7F9C3),
   .weight25_2_pe0(24'h5E2F07),
   .weight26_2_pe0(24'h7F1027),
   .weight27_2_pe0(24'h3113E5),
   .weight28_2_pe0(24'h808080),
   .weight29_2_pe0(24'h808080),
   .weight30_2_pe0(24'h808080),
   .weight31_2_pe0(24'hA4300F),
   .weight32_2_pe0(24'hEC18F5),
   .weight33_2_pe0(24'hDFEBE2),
   .weight34_2_pe0(24'h170E1F),
   .weight35_2_pe0(24'hE51830),
   .weight36_2_pe0(24'hFE811C),
   .weight01_1_pe1(24'h2BFF2A),
   .weight02_1_pe1(24'h11CA16),
   .weight03_1_pe1(24'hEDD4EE),
   .weight04_1_pe1(24'h279FC0),
   .weight05_1_pe1(24'h001DA3),
   .weight06_1_pe1(24'h1B2B0E),
   .weight07_1_pe1(24'hCB2AED),
   .weight08_1_pe1(24'hF20BE4),
   .weight09_1_pe1(24'h2815FB),
   .weight10_1_pe1(24'h0CF6D2),
   .weight11_1_pe1(24'hD97FD8),
   .weight12_1_pe1(24'hF5E0D9),
   .weight13_1_pe1(24'h11F8F0),
   .weight14_1_pe1(24'h126D1C),
   .weight15_1_pe1(24'h1BF709),
   .weight16_1_pe1(24'h0E0A0B),
   .weight17_1_pe1(24'hD7FC05),
   .weight18_1_pe1(24'h14FA11),
   .weight19_1_pe1(24'hC4BE0A),
   .weight20_1_pe1(24'hD29211),
   .weight21_1_pe1(24'hF3072B),
   .weight22_1_pe1(24'h1FCBFD),
   .weight23_1_pe1(24'hFB7F18),
   .weight24_1_pe1(24'h1616F8),
   .weight25_1_pe1(24'hF24309),
   .weight26_1_pe1(24'hE728D3),
   .weight27_1_pe1(24'h110604),
   .weight28_1_pe1(24'h17FDDB),
   .weight29_1_pe1(24'h01F21F),
   .weight30_1_pe1(24'hF10E17),
   .weight31_1_pe1(24'hD8220D),
   .weight32_1_pe1(24'h0B2F14),
   .weight33_1_pe1(24'hF1EDF1),
   .weight34_1_pe1(24'hFC26F5),
   .weight35_1_pe1(24'hF85EFB),
   .weight36_1_pe1(24'hE6F4F0),
   .weight01_2_pe1(24'h52E6DA),
   .weight02_2_pe1(24'h572ACC),
   .weight03_2_pe1(24'h2079C8),
   .weight04_2_pe1(24'h80007F),
   .weight05_2_pe1(24'h8019BE),
   .weight06_2_pe1(24'hFCB706),
   .weight07_2_pe1(24'hE305E1),
   .weight08_2_pe1(24'hE92608),
   .weight09_2_pe1(24'hC0E903),
   .weight10_2_pe1(24'hAEE71F),
   .weight11_2_pe1(24'h2F7E1B),
   .weight12_2_pe1(24'h2DE68D),
   .weight13_2_pe1(24'h9BF3D3),
   .weight14_2_pe1(24'hC97E01),
   .weight15_2_pe1(24'hD6DEB2),
   .weight16_2_pe1(24'h2B12E8),
   .weight17_2_pe1(24'hD87FB7),
   .weight18_2_pe1(24'hFB4D7F),
   .weight19_2_pe1(24'h6EF5FA),
   .weight20_2_pe1(24'h0980E2),
   .weight21_2_pe1(24'h190DE0),
   .weight22_2_pe1(24'hE99DEC),
   .weight23_2_pe1(24'h1E0945),
   .weight24_2_pe1(24'h04E320),
   .weight25_2_pe1(24'hE742F4),
   .weight26_2_pe1(24'hCEBEC6),
   .weight27_2_pe1(24'hF6292F),
   .weight28_2_pe1(24'h00F87F),
   .weight29_2_pe1(24'h7E7F6E),
   .weight30_2_pe1(24'h1EDD80),
   .weight31_2_pe1(24'h7F561D),
   .weight32_2_pe1(24'hC7F207),
   .weight33_2_pe1(24'h1C1CFF),
   .weight34_2_pe1(24'hDD59DF),
   .weight35_2_pe1(24'h210153),
   .weight36_2_pe1(24'h21D708),
   .weight01_1_pe2(24'hC135DA),
   .weight02_1_pe2(24'h802AD2),
   .weight03_1_pe2(24'h2F41F0),
   .weight04_1_pe2(24'h7FBD4D),
   .weight05_1_pe2(24'h04E920),
   .weight06_1_pe2(24'hCCCBF6),
   .weight07_1_pe2(24'hEBF10E),
   .weight08_1_pe2(24'hDD36F2),
   .weight09_1_pe2(24'hE9EC24),
   .weight10_1_pe2(24'h0EF2F9),
   .weight11_1_pe2(24'h0A5AEF),
   .weight12_1_pe2(24'h2D0C0E),
   .weight13_1_pe2(24'h0E4CEF),
   .weight14_1_pe2(24'h134F2D),
   .weight15_1_pe2(24'hF6B91D),
   .weight16_1_pe2(24'h0607D8),
   .weight17_1_pe2(24'hBB570B),
   .weight18_1_pe2(24'hF6D7E9),
   .weight19_1_pe2(24'h2DF319),
   .weight20_1_pe2(24'hE97F12),
   .weight21_1_pe2(24'hEAD9CC),
   .weight22_1_pe2(24'h201622),
   .weight23_1_pe2(24'h0556F3),
   .weight24_1_pe2(24'hE1FDEA),
   .weight25_1_pe2(24'hFD03E8),
   .weight26_1_pe2(24'hF75B1A),
   .weight27_1_pe2(24'hF225F8),
   .weight28_1_pe2(24'h21190B),
   .weight29_1_pe2(24'hFD80A5),
   .weight30_1_pe2(24'hF71C2A),
   .weight31_1_pe2(24'hF7E1ED),
   .weight32_1_pe2(24'h1439BD),
   .weight33_1_pe2(24'h0F07F1),
   .weight34_1_pe2(24'hF4F2F6),
   .weight35_1_pe2(24'hDC540D),
   .weight36_1_pe2(24'h1BDD02),
   .weight01_2_pe2(24'hF6CB64),
   .weight02_2_pe2(24'h38F5BE),
   .weight03_2_pe2(24'hDECE24),
   .weight04_2_pe2(24'h808291),
   .weight05_2_pe2(24'hDB6228),
   .weight06_2_pe2(24'h4B06E6),
   .weight07_2_pe2(24'h2E12D2),
   .weight08_2_pe2(24'h0F5FE6),
   .weight09_2_pe2(24'h4026FF),
   .weight10_2_pe2(24'h0413FD),
   .weight11_2_pe2(24'h1A70BD),
   .weight12_2_pe2(24'hFA13E2),
   .weight13_2_pe2(24'hEC34DB),
   .weight14_2_pe2(24'h2025ED),
   .weight15_2_pe2(24'h014FF6),
   .weight16_2_pe2(24'hC7D717),
   .weight17_2_pe2(24'h0A3E27),
   .weight18_2_pe2(24'hFCE860),
   .weight19_2_pe2(24'h043CF1),
   .weight20_2_pe2(24'hF3D0ED),
   .weight21_2_pe2(24'h7FC1D3),
   .weight22_2_pe2(24'h12E4FE),
   .weight23_2_pe2(24'hFB01F9),
   .weight24_2_pe2(24'h1526AE),
   .weight25_2_pe2(24'hD125C7),
   .weight26_2_pe2(24'h45F112),
   .weight27_2_pe2(24'hE90609),
   .weight28_2_pe2(24'hF5E9D7),
   .weight29_2_pe2(24'h31270B),
   .weight30_2_pe2(24'h0C1E82),
   .weight31_2_pe2(24'hE90818),
   .weight32_2_pe2(24'hF8250D),
   .weight33_2_pe2(24'h040508),
   .weight34_2_pe2(24'h380115),
   .weight35_2_pe2(24'h3CCE52),
   .weight36_2_pe2(24'h900906),
   .weight01_1_pe3(24'h80BCFE),
   .weight02_1_pe3(24'h7F7FB3),
   .weight03_1_pe3(24'hEBC11C),
   .weight04_1_pe3(24'h547F78),
   .weight05_1_pe3(24'h808080),
   .weight06_1_pe3(24'hD47F80),
   .weight07_1_pe3(24'h2E7F1E),
   .weight08_1_pe3(24'h1A8082),
   .weight09_1_pe3(24'h807F7F),
   .weight10_1_pe3(24'h0B79E7),
   .weight11_1_pe3(24'h357FB6),
   .weight12_1_pe3(24'h5B8031),
   .weight13_1_pe3(24'hC4CB80),
   .weight14_1_pe3(24'h2B583D),
   .weight15_1_pe3(24'h11800F),
   .weight16_1_pe3(24'hF91904),
   .weight17_1_pe3(24'hF27F7F),
   .weight18_1_pe3(24'h0E807F),
   .weight19_1_pe3(24'h6E7F62),
   .weight20_1_pe3(24'hCC51EA),
   .weight21_1_pe3(24'h8F8080),
   .weight22_1_pe3(24'h1CAF7F),
   .weight23_1_pe3(24'hAC7E2A),
   .weight24_1_pe3(24'hBF040E),
   .weight25_1_pe3(24'h507EBE),
   .weight26_1_pe3(24'h54BE35),
   .weight27_1_pe3(24'hAB1CF8),
   .weight28_1_pe3(24'hFE7644),
   .weight29_1_pe3(24'h2CD59E),
   .weight30_1_pe3(24'h6D7D76),
   .weight31_1_pe3(24'h037E88),
   .weight32_1_pe3(24'hE280CB),
   .weight33_1_pe3(24'hF70B80),
   .weight34_1_pe3(24'hE780AC),
   .weight35_1_pe3(24'h807F5E),
   .weight36_1_pe3(24'h7F80B2),
   .weight01_2_pe3(24'h108041),
   .weight02_2_pe3(24'h107F21),
   .weight03_2_pe3(24'h110804),
   .weight04_2_pe3(24'hABC3A4),
   .weight05_2_pe3(24'hD3BBE9),
   .weight06_2_pe3(24'hFB1ED5),
   .weight07_2_pe3(24'hD346DC),
   .weight08_2_pe3(24'hAE7F27),
   .weight09_2_pe3(24'hADB87F),
   .weight10_2_pe3(24'hFBE60E),
   .weight11_2_pe3(24'h053FF6),
   .weight12_2_pe3(24'h17F5F0),
   .weight13_2_pe3(24'hA513DA),
   .weight14_2_pe3(24'hD324EE),
   .weight15_2_pe3(24'hCA09ED),
   .weight16_2_pe3(24'hFC1FF8),
   .weight17_2_pe3(24'h0335FB),
   .weight18_2_pe3(24'h04AF64),
   .weight19_2_pe3(24'hBEE914),
   .weight20_2_pe3(24'h120C25),
   .weight21_2_pe3(24'h019DCB),
   .weight22_2_pe3(24'hBFDBED),
   .weight23_2_pe3(24'hDF7431),
   .weight24_2_pe3(24'hD9BA56),
   .weight25_2_pe3(24'h3F09DF),
   .weight26_2_pe3(24'h4EDD25),
   .weight27_2_pe3(24'hFAFBE9),
   .weight28_2_pe3(24'hE1FE05),
   .weight29_2_pe3(24'hEB11D9),
   .weight30_2_pe3(24'h277F0D),
   .weight31_2_pe3(24'h4737D1),
   .weight32_2_pe3(24'h6526CB),
   .weight33_2_pe3(24'h1341DF),
   .weight34_2_pe3(24'h59F91F),
   .weight35_2_pe3(24'hEA0631),
   .weight36_2_pe3(24'h0CE11B),
   .weight01_1_pe4(24'hD561AD),
   .weight02_1_pe4(24'hE39151),
   .weight03_1_pe4(24'hF91136),
   .weight04_1_pe4(24'h7F7F7F),
   .weight05_1_pe4(24'h617F77),
   .weight06_1_pe4(24'hF0FC06),
   .weight07_1_pe4(24'h1DD2F0),
   .weight08_1_pe4(24'h398036),
   .weight09_1_pe4(24'h02AEE0),
   .weight10_1_pe4(24'hE1AB2B),
   .weight11_1_pe4(24'hE63122),
   .weight12_1_pe4(24'h4BFC5F),
   .weight13_1_pe4(24'h22F5FD),
   .weight14_1_pe4(24'hC97FF9),
   .weight15_1_pe4(24'hF023F0),
   .weight16_1_pe4(24'h0FE52B),
   .weight17_1_pe4(24'h1BF5DC),
   .weight18_1_pe4(24'h0AA1CB),
   .weight19_1_pe4(24'hAE150C),
   .weight20_1_pe4(24'h80F4F7),
   .weight21_1_pe4(24'hEA43FA),
   .weight22_1_pe4(24'hC4F4D4),
   .weight23_1_pe4(24'h1EF71A),
   .weight24_1_pe4(24'hFFF225),
   .weight25_1_pe4(24'h20977F),
   .weight26_1_pe4(24'h7FB8D1),
   .weight27_1_pe4(24'h2FDDE2),
   .weight28_1_pe4(24'hE72508),
   .weight29_1_pe4(24'hFD147F),
   .weight30_1_pe4(24'hF0E77F),
   .weight31_1_pe4(24'hF87603),
   .weight32_1_pe4(24'hCD4131),
   .weight33_1_pe4(24'h072F11),
   .weight34_1_pe4(24'hEB0ADA),
   .weight35_1_pe4(24'hEE34D0),
   .weight36_1_pe4(24'h081E01),
   .weight01_2_pe4(24'hE953F1),
   .weight02_2_pe4(24'h7F7FEF),
   .weight03_2_pe4(24'h5BCB23),
   .weight04_2_pe4(24'hEDA3C8),
   .weight05_2_pe4(24'hED8162),
   .weight06_2_pe4(24'hB17B04),
   .weight07_2_pe4(24'h6D7F03),
   .weight08_2_pe4(24'h7FDE03),
   .weight09_2_pe4(24'hDA7FEA),
   .weight10_2_pe4(24'hDE1032),
   .weight11_2_pe4(24'hCC7F03),
   .weight12_2_pe4(24'h837069),
   .weight13_2_pe4(24'h09ADC3),
   .weight14_2_pe4(24'hCCBB43),
   .weight15_2_pe4(24'hFE12F4),
   .weight16_2_pe4(24'h2A2BF4),
   .weight17_2_pe4(24'h37E615),
   .weight18_2_pe4(24'h255E14),
   .weight19_2_pe4(24'hF8043C),
   .weight20_2_pe4(24'h655C02),
   .weight21_2_pe4(24'h8D4BE8),
   .weight22_2_pe4(24'h31830A),
   .weight23_2_pe4(24'h257FD5),
   .weight24_2_pe4(24'hA37782),
   .weight25_2_pe4(24'hDCE9F8),
   .weight26_2_pe4(24'h748150),
   .weight27_2_pe4(24'h060EC5),
   .weight28_2_pe4(24'hEE28DD),
   .weight29_2_pe4(24'hA60B74),
   .weight30_2_pe4(24'h1B167F),
   .weight31_2_pe4(24'h167FF2),
   .weight32_2_pe4(24'h108024),
   .weight33_2_pe4(24'h1AF518),
   .weight34_2_pe4(24'h25F10C),
   .weight35_2_pe4(24'h82D9D4),
   .weight36_2_pe4(24'h17AB0F),
   .weight01_1_pe5(24'h44BDEE),
   .weight02_1_pe5(24'hC75609),
   .weight03_1_pe5(24'hF1FAFD),
   .weight04_1_pe5(24'h497FEA),
   .weight05_1_pe5(24'h2CE9C4),
   .weight06_1_pe5(24'hE50718),
   .weight07_1_pe5(24'hF91335),
   .weight08_1_pe5(24'hDA9B0C),
   .weight09_1_pe5(24'h1305DE),
   .weight10_1_pe5(24'hD72019),
   .weight11_1_pe5(24'hE67EC5),
   .weight12_1_pe5(24'hF205D1),
   .weight13_1_pe5(24'hCFE3F0),
   .weight14_1_pe5(24'hE65BD0),
   .weight15_1_pe5(24'hF307EE),
   .weight16_1_pe5(24'h2A3322),
   .weight17_1_pe5(24'hD52B16),
   .weight18_1_pe5(24'h0F0A06),
   .weight19_1_pe5(24'h7F3CDF),
   .weight20_1_pe5(24'h7F2604),
   .weight21_1_pe5(24'h222E51),
   .weight22_1_pe5(24'hEBF41D),
   .weight23_1_pe5(24'h062515),
   .weight24_1_pe5(24'h1F07EF),
   .weight25_1_pe5(24'h383BE6),
   .weight26_1_pe5(24'h183B26),
   .weight27_1_pe5(24'hF3060A),
   .weight28_1_pe5(24'hF3F7F5),
   .weight29_1_pe5(24'h04EDE6),
   .weight30_1_pe5(24'hFEE880),
   .weight31_1_pe5(24'h17D406),
   .weight32_1_pe5(24'h083C12),
   .weight33_1_pe5(24'hF8CF09),
   .weight34_1_pe5(24'hF7F21C),
   .weight35_1_pe5(24'hC743F0),
   .weight36_1_pe5(24'h34F417),
   .weight01_2_pe5(24'h2616DA),
   .weight02_2_pe5(24'h7F800D),
   .weight03_2_pe5(24'h64EBF2),
   .weight04_2_pe5(24'h29F0F9),
   .weight05_2_pe5(24'h7F78EF),
   .weight06_2_pe5(24'h80FEF4),
   .weight07_2_pe5(24'hFDBFF9),
   .weight08_2_pe5(24'h7F070E),
   .weight09_2_pe5(24'h9F0300),
   .weight10_2_pe5(24'hEAB920),
   .weight11_2_pe5(24'h817F80),
   .weight12_2_pe5(24'h80370F),
   .weight13_2_pe5(24'hBB7FA5),
   .weight14_2_pe5(24'h80D363),
   .weight15_2_pe5(24'h80FA80),
   .weight16_2_pe5(24'h0AFCDB),
   .weight17_2_pe5(24'hAC7F1F),
   .weight18_2_pe5(24'h808009),
   .weight19_2_pe5(24'h98FBF4),
   .weight20_2_pe5(24'h8080FB),
   .weight21_2_pe5(24'h7F80EF),
   .weight22_2_pe5(24'h7FD21D),
   .weight23_2_pe5(24'h1D285D),
   .weight24_2_pe5(24'h8262C3),
   .weight25_2_pe5(24'h801403),
   .weight26_2_pe5(24'h80C60A),
   .weight27_2_pe5(24'h807FCC),
   .weight28_2_pe5(24'h2C080E),
   .weight29_2_pe5(24'h437FE1),
   .weight30_2_pe5(24'h8080F5),
   .weight31_2_pe5(24'hC46BE3),
   .weight32_2_pe5(24'h823AFB),
   .weight33_2_pe5(24'h7BE751),
   .weight34_2_pe5(24'hDB361C),
   .weight35_2_pe5(24'h7F7F35),
   .weight36_2_pe5(24'h7F9200)
)core_layer1(
   .i_clk(i_clk),
   .i_rstn(i_rstn),
   .s_axis_tready(s_axis_tready),
   .s_axis_tvalid(s_axis_tvalid),
   .s_axis_tdata(s_axis_tdata),
   .m_axis_tdata(m_axis_tdata_core[0]),
   .m_axis_tvalid(m_axis_tvalid_core[0]),
   .m_axis_tready(m_axis_tready_core[0]),
   .EOL(),
   .EOF()
);

Axi4ConvCore#(
   .REQUANT(77),
   .weight01_1_pe0(24'hC557CF),
   .weight02_1_pe0(24'hFF09D9),
   .weight03_1_pe0(24'h387E07),
   .weight04_1_pe0(24'h7F5D83),
   .weight05_1_pe0(24'h668080),
   .weight06_1_pe0(24'h6E7FF3),
   .weight07_1_pe0(24'hC1C8FA),
   .weight08_1_pe0(24'h807FB5),
   .weight09_1_pe0(24'h80BC16),
   .weight10_1_pe0(24'hA75030),
   .weight11_1_pe0(24'h808068),
   .weight12_1_pe0(24'hF4F3CC),
   .weight13_1_pe0(24'h09AE31),
   .weight14_1_pe0(24'h7FF462),
   .weight15_1_pe0(24'hCC3E91),
   .weight16_1_pe0(24'hCA077F),
   .weight17_1_pe0(24'h0C816C),
   .weight18_1_pe0(24'h80ABDF),
   .weight19_1_pe0(24'hEFADAD),
   .weight20_1_pe0(24'hC1B9E0),
   .weight21_1_pe0(24'h807207),
   .weight22_1_pe0(24'h70FA40),
   .weight23_1_pe0(24'h7F8032),
   .weight24_1_pe0(24'h7B7FF8),
   .weight25_1_pe0(24'hF8B086),
   .weight26_1_pe0(24'hE7CDC4),
   .weight27_1_pe0(24'h617F1F),
   .weight28_1_pe0(24'hF1A665),
   .weight29_1_pe0(24'hD5B857),
   .weight30_1_pe0(24'h497F7F),
   .weight31_1_pe0(24'h2F7F07),
   .weight32_1_pe0(24'h99804C),
   .weight33_1_pe0(24'h7F7F5A),
   .weight34_1_pe0(24'hA532F9),
   .weight35_1_pe0(24'hFE0C7F),
   .weight36_1_pe0(24'h04FCB9),
   .weight01_2_pe0(24'h2CFB23),
   .weight02_2_pe0(24'h1C1C12),
   .weight03_2_pe0(24'h020C59),
   .weight04_2_pe0(24'hD808AF),
   .weight05_2_pe0(24'h177F2B),
   .weight06_2_pe0(24'hEE612E),
   .weight07_2_pe0(24'h0E5919),
   .weight08_2_pe0(24'hDE7F36),
   .weight09_2_pe0(24'h870F9F),
   .weight10_2_pe0(24'h28DE49),
   .weight11_2_pe0(24'h9A05D2),
   .weight12_2_pe0(24'h249C10),
   .weight13_2_pe0(24'h286168),
   .weight14_2_pe0(24'h0C281D),
   .weight15_2_pe0(24'h978009),
   .weight16_2_pe0(24'hB67F13),
   .weight17_2_pe0(24'hE57FEA),
   .weight18_2_pe0(24'h0D8022),
   .weight19_2_pe0(24'h1580F4),
   .weight20_2_pe0(24'h7FB241),
   .weight21_2_pe0(24'h3DF12D),
   .weight22_2_pe0(24'hEA2F25),
   .weight23_2_pe0(24'hE27EF8),
   .weight24_2_pe0(24'hB8B91A),
   .weight25_2_pe0(24'hCDF1B7),
   .weight26_2_pe0(24'h167FC9),
   .weight27_2_pe0(24'h0B101C),
   .weight28_2_pe0(24'h29CA90),
   .weight29_2_pe0(24'h1F7F00),
   .weight30_2_pe0(24'h054818),
   .weight31_2_pe0(24'hCEBB6A),
   .weight32_2_pe0(24'hF04CB9),
   .weight33_2_pe0(24'hEBF71F),
   .weight34_2_pe0(24'h1F807F),
   .weight35_2_pe0(24'h05E35D),
   .weight36_2_pe0(24'hEBF8FD),
   .weight01_1_pe1(24'hE6F807),
   .weight02_1_pe1(24'hE70CE5),
   .weight03_1_pe1(24'hF5F008),
   .weight04_1_pe1(24'hEFF8FF),
   .weight05_1_pe1(24'hEEF7FA),
   .weight06_1_pe1(24'hFA01DF),
   .weight07_1_pe1(24'hFCF8F5),
   .weight08_1_pe1(24'h1812EB),
   .weight09_1_pe1(24'hF801F5),
   .weight10_1_pe1(24'h1A020C),
   .weight11_1_pe1(24'hF0FD10),
   .weight12_1_pe1(24'hF407F0),
   .weight13_1_pe1(24'hF2EB07),
   .weight14_1_pe1(24'hF903FD),
   .weight15_1_pe1(24'hF10EFE),
   .weight16_1_pe1(24'hE814FA),
   .weight17_1_pe1(24'hFBF0F4),
   .weight18_1_pe1(24'h0306FC),
   .weight19_1_pe1(24'h0CF2E1),
   .weight20_1_pe1(24'hF0FDFE),
   .weight21_1_pe1(24'h19F214),
   .weight22_1_pe1(24'h05EE06),
   .weight23_1_pe1(24'hF4EDF0),
   .weight24_1_pe1(24'hFCEFEE),
   .weight25_1_pe1(24'hF80DF3),
   .weight26_1_pe1(24'h020608),
   .weight27_1_pe1(24'hF614EF),
   .weight28_1_pe1(24'h0CF6F7),
   .weight29_1_pe1(24'hECED03),
   .weight30_1_pe1(24'hFCE703),
   .weight31_1_pe1(24'hED04F5),
   .weight32_1_pe1(24'h14F5ED),
   .weight33_1_pe1(24'h02EF13),
   .weight34_1_pe1(24'h0BEF04),
   .weight35_1_pe1(24'hE5EDFC),
   .weight36_1_pe1(24'hF1E5E3),
   .weight01_2_pe1(24'h44A111),
   .weight02_2_pe1(24'hE406D0),
   .weight03_2_pe1(24'h22BDE7),
   .weight04_2_pe1(24'hE1E032),
   .weight05_2_pe1(24'h237F16),
   .weight06_2_pe1(24'hF704F4),
   .weight07_2_pe1(24'hE9EA0A),
   .weight08_2_pe1(24'h0D7F3C),
   .weight09_2_pe1(24'h64320B),
   .weight10_2_pe1(24'hD45CD9),
   .weight11_2_pe1(24'h7FA4FC),
   .weight12_2_pe1(24'hB01202),
   .weight13_2_pe1(24'h1536E8),
   .weight14_2_pe1(24'hD27F45),
   .weight15_2_pe1(24'h2B030B),
   .weight16_2_pe1(24'hCF1CFA),
   .weight17_2_pe1(24'h236D2E),
   .weight18_2_pe1(24'hF7440F),
   .weight19_2_pe1(24'h2D1EEC),
   .weight20_2_pe1(24'hFB7F1C),
   .weight21_2_pe1(24'hDA9B0B),
   .weight22_2_pe1(24'hEAEA41),
   .weight23_2_pe1(24'hEA44EE),
   .weight24_2_pe1(24'h0FFF06),
   .weight25_2_pe1(24'h04E601),
   .weight26_2_pe1(24'h2875FE),
   .weight27_2_pe1(24'hD2BE9A),
   .weight28_2_pe1(24'hEEB103),
   .weight29_2_pe1(24'hD048BC),
   .weight30_2_pe1(24'h20E3E1),
   .weight31_2_pe1(24'h1D0D53),
   .weight32_2_pe1(24'hE77FB3),
   .weight33_2_pe1(24'hFD17F5),
   .weight34_2_pe1(24'h3BF880),
   .weight35_2_pe1(24'hD74280),
   .weight36_2_pe1(24'hF41F0E),
   .weight01_1_pe2(24'h8E0436),
   .weight02_1_pe2(24'h3B7F35),
   .weight03_1_pe2(24'hD418F5),
   .weight04_1_pe2(24'h7F3B22),
   .weight05_1_pe2(24'h3A7089),
   .weight06_1_pe2(24'h90C116),
   .weight07_1_pe2(24'h126E24),
   .weight08_1_pe2(24'h7F7FB5),
   .weight09_1_pe2(24'h7C9FA4),
   .weight10_1_pe2(24'h0F3BEC),
   .weight11_1_pe2(24'h688228),
   .weight12_1_pe2(24'hFA3C02),
   .weight13_1_pe2(24'hC2809C),
   .weight14_1_pe2(24'h9F80D8),
   .weight15_1_pe2(24'h40B226),
   .weight16_1_pe2(24'h996345),
   .weight17_1_pe2(24'hD0A504),
   .weight18_1_pe2(24'h02F43B),
   .weight19_1_pe2(24'h7FAF26),
   .weight20_1_pe2(24'h7F9822),
   .weight21_1_pe2(24'h4AD266),
   .weight22_1_pe2(24'h7F25E3),
   .weight23_1_pe2(24'h2D9059),
   .weight24_1_pe2(24'hEF1CE9),
   .weight25_1_pe2(24'h90808F),
   .weight26_1_pe2(24'h7FCA00),
   .weight27_1_pe2(24'h3762DF),
   .weight28_1_pe2(24'hD17F38),
   .weight29_1_pe2(24'h7F8199),
   .weight30_1_pe2(24'hA9A574),
   .weight31_1_pe2(24'h5D7F09),
   .weight32_1_pe2(24'hCD807F),
   .weight33_1_pe2(24'hE26259),
   .weight34_1_pe2(24'hC27F7F),
   .weight35_1_pe2(24'h00387F),
   .weight36_1_pe2(24'hE621B8),
   .weight01_2_pe2(24'h31F900),
   .weight02_2_pe2(24'hE2650B),
   .weight03_2_pe2(24'h0EEE26),
   .weight04_2_pe2(24'hEFFDE8),
   .weight05_2_pe2(24'h437F30),
   .weight06_2_pe2(24'h20F0CF),
   .weight07_2_pe2(24'h2E3D03),
   .weight08_2_pe2(24'h147FC2),
   .weight09_2_pe2(24'h00F701),
   .weight10_2_pe2(24'hD727B3),
   .weight11_2_pe2(24'h2F0913),
   .weight12_2_pe2(24'h23E8F2),
   .weight13_2_pe2(24'hFA4F95),
   .weight14_2_pe2(24'hCB7FDD),
   .weight15_2_pe2(24'h0AD2F6),
   .weight16_2_pe2(24'h351CD6),
   .weight17_2_pe2(24'h107F0E),
   .weight18_2_pe2(24'h2CF9F2),
   .weight19_2_pe2(24'h97C54A),
   .weight20_2_pe2(24'hA5B27D),
   .weight21_2_pe2(24'h1D56EF),
   .weight22_2_pe2(24'hE5191A),
   .weight23_2_pe2(24'hB67202),
   .weight24_2_pe2(24'h102075),
   .weight25_2_pe2(24'h22E53C),
   .weight26_2_pe2(24'h367615),
   .weight27_2_pe2(24'h142418),
   .weight28_2_pe2(24'hB7C0F7),
   .weight29_2_pe2(24'h846CCC),
   .weight30_2_pe2(24'hD106C7),
   .weight31_2_pe2(24'hE5C532),
   .weight32_2_pe2(24'hFE5CE5),
   .weight33_2_pe2(24'hFCE6D3),
   .weight34_2_pe2(24'hF48080),
   .weight35_2_pe2(24'h095010),
   .weight36_2_pe2(24'hD5D8B6),
   .weight01_1_pe3(24'hABCFFB),
   .weight02_1_pe3(24'h53AD15),
   .weight03_1_pe3(24'hF336E2),
   .weight04_1_pe3(24'h7F7F51),
   .weight05_1_pe3(24'hC88372),
   .weight06_1_pe3(24'h7F3D1A),
   .weight07_1_pe3(24'hCD7F80),
   .weight08_1_pe3(24'h8FB0EA),
   .weight09_1_pe3(24'hC531A2),
   .weight10_1_pe3(24'hE84F23),
   .weight11_1_pe3(24'h153DBC),
   .weight12_1_pe3(24'h2A4142),
   .weight13_1_pe3(24'h555D0D),
   .weight14_1_pe3(24'h7F617F),
   .weight15_1_pe3(24'h145B3C),
   .weight16_1_pe3(24'h808380),
   .weight17_1_pe3(24'h828198),
   .weight18_1_pe3(24'hDEB71D),
   .weight19_1_pe3(24'h808080),
   .weight20_1_pe3(24'h068080),
   .weight21_1_pe3(24'h95A0D2),
   .weight22_1_pe3(24'h7D79F1),
   .weight23_1_pe3(24'h03857F),
   .weight24_1_pe3(24'h0C7FE4),
   .weight25_1_pe3(24'h04ED1C),
   .weight26_1_pe3(24'h108010),
   .weight27_1_pe3(24'hB6B534),
   .weight28_1_pe3(24'h2A7F80),
   .weight29_1_pe3(24'h024F7F),
   .weight30_1_pe3(24'h7F80FF),
   .weight31_1_pe3(24'h182897),
   .weight32_1_pe3(24'h21817F),
   .weight33_1_pe3(24'hCFBCDA),
   .weight34_1_pe3(24'h072F7F),
   .weight35_1_pe3(24'h26427E),
   .weight36_1_pe3(24'hFDF3FA),
   .weight01_2_pe3(24'hD280D8),
   .weight02_2_pe3(24'h8080C5),
   .weight03_2_pe3(24'hD3801B),
   .weight04_2_pe3(24'h4D005C),
   .weight05_2_pe3(24'h5E7F30),
   .weight06_2_pe3(24'h4B7F00),
   .weight07_2_pe3(24'hE980C2),
   .weight08_2_pe3(24'h7B7F7F),
   .weight09_2_pe3(24'h287F41),
   .weight10_2_pe3(24'hF706EF),
   .weight11_2_pe3(24'h146202),
   .weight12_2_pe3(24'h161A3B),
   .weight13_2_pe3(24'h0B7F1A),
   .weight14_2_pe3(24'hFA7F5C),
   .weight15_2_pe3(24'h2FEE0A),
   .weight16_2_pe3(24'hD1F781),
   .weight17_2_pe3(24'h8C7FDE),
   .weight18_2_pe3(24'h3E18D2),
   .weight19_2_pe3(24'h3B1DF0),
   .weight20_2_pe3(24'h7F7F0B),
   .weight21_2_pe3(24'hB641DC),
   .weight22_2_pe3(24'h2BC2E2),
   .weight23_2_pe3(24'h4E7FD3),
   .weight24_2_pe3(24'hFD892A),
   .weight25_2_pe3(24'h084F75),
   .weight26_2_pe3(24'hCB7F2B),
   .weight27_2_pe3(24'hDA26F5),
   .weight28_2_pe3(24'h474714),
   .weight29_2_pe3(24'hA27FEB),
   .weight30_2_pe3(24'hDF8884),
   .weight31_2_pe3(24'h8980A1),
   .weight32_2_pe3(24'hF57F80),
   .weight33_2_pe3(24'hEA809F),
   .weight34_2_pe3(24'hFD4D50),
   .weight35_2_pe3(24'h2B7F89),
   .weight36_2_pe3(24'h171033),
   .weight01_1_pe4(24'hED25D4),
   .weight02_1_pe4(24'h064531),
   .weight03_1_pe4(24'hEDDA03),
   .weight04_1_pe4(24'hF3DEED),
   .weight05_1_pe4(24'hEB7F5C),
   .weight06_1_pe4(24'hD9DCD8),
   .weight07_1_pe4(24'h3708FB),
   .weight08_1_pe4(24'h0D7F60),
   .weight09_1_pe4(24'h3EE701),
   .weight10_1_pe4(24'hC8FC1D),
   .weight11_1_pe4(24'hE652E9),
   .weight12_1_pe4(24'hE909FB),
   .weight13_1_pe4(24'hEB2B0F),
   .weight14_1_pe4(24'hD57D13),
   .weight15_1_pe4(24'hE6F7E4),
   .weight16_1_pe4(24'hE2E7ED),
   .weight17_1_pe4(24'hFF7F22),
   .weight18_1_pe4(24'hEB07E0),
   .weight19_1_pe4(24'hB55BCD),
   .weight20_1_pe4(24'h1CE0D4),
   .weight21_1_pe4(24'hE8E0E6),
   .weight22_1_pe4(24'h27D5DA),
   .weight23_1_pe4(24'h0838D5),
   .weight24_1_pe4(24'h42CBE7),
   .weight25_1_pe4(24'hE713D4),
   .weight26_1_pe4(24'hAF7FCA),
   .weight27_1_pe4(24'hC40AFD),
   .weight28_1_pe4(24'h1F12E6),
   .weight29_1_pe4(24'hEB7722),
   .weight30_1_pe4(24'h463B22),
   .weight31_1_pe4(24'h47D9F1),
   .weight32_1_pe4(24'h3175FD),
   .weight33_1_pe4(24'hEC25D4),
   .weight34_1_pe4(24'h33EB7F),
   .weight35_1_pe4(24'h01BBFA),
   .weight36_1_pe4(24'h13C257),
   .weight01_2_pe4(24'hE62312),
   .weight02_2_pe4(24'hAB2BD5),
   .weight03_2_pe4(24'h36CFFE),
   .weight04_2_pe4(24'h2D1E0F),
   .weight05_2_pe4(24'hEC7F2F),
   .weight06_2_pe4(24'hF0300B),
   .weight07_2_pe4(24'hE70ED7),
   .weight08_2_pe4(24'h257F60),
   .weight09_2_pe4(24'hFFD4FC),
   .weight10_2_pe4(24'h344019),
   .weight11_2_pe4(24'hE68107),
   .weight12_2_pe4(24'h11410D),
   .weight13_2_pe4(24'hFCF3F2),
   .weight14_2_pe4(24'hD37F00),
   .weight15_2_pe4(24'h23E30C),
   .weight16_2_pe4(24'h11F0ED),
   .weight17_2_pe4(24'hFA7F15),
   .weight18_2_pe4(24'hF156DB),
   .weight19_2_pe4(24'hEBF52A),
   .weight20_2_pe4(24'hB94CCE),
   .weight21_2_pe4(24'h56BD3D),
   .weight22_2_pe4(24'hFDE0F5),
   .weight23_2_pe4(24'h017D0A),
   .weight24_2_pe4(24'h16DACD),
   .weight25_2_pe4(24'hD71D0A),
   .weight26_2_pe4(24'h2A7FF8),
   .weight27_2_pe4(24'hCFE2FB),
   .weight28_2_pe4(24'hFDF224),
   .weight29_2_pe4(24'h237A20),
   .weight30_2_pe4(24'hE7F5E9),
   .weight31_2_pe4(24'hFCC1E0),
   .weight32_2_pe4(24'h087FF7),
   .weight33_2_pe4(24'hF8D5C6),
   .weight34_2_pe4(24'hDCC7AA),
   .weight35_2_pe4(24'hF74E80),
   .weight36_2_pe4(24'hEFDD45),
   .weight01_1_pe5(24'hF514DE),
   .weight02_1_pe5(24'hBDC2D8),
   .weight03_1_pe5(24'h2C0929),
   .weight04_1_pe5(24'h25EADE),
   .weight05_1_pe5(24'h5C7F2A),
   .weight06_1_pe5(24'h1C43F8),
   .weight07_1_pe5(24'hDD16C8),
   .weight08_1_pe5(24'hF67C04),
   .weight09_1_pe5(24'hD90E10),
   .weight10_1_pe5(24'hE3A21B),
   .weight11_1_pe5(24'h190B1C),
   .weight12_1_pe5(24'h05EDF9),
   .weight13_1_pe5(24'hEDAFF2),
   .weight14_1_pe5(24'hF47FE0),
   .weight15_1_pe5(24'hEF0A05),
   .weight16_1_pe5(24'hD2E40D),
   .weight17_1_pe5(24'h2878F9),
   .weight18_1_pe5(24'hE406CD),
   .weight19_1_pe5(24'h470BDF),
   .weight20_1_pe5(24'h12C4C5),
   .weight21_1_pe5(24'hB723E3),
   .weight22_1_pe5(24'h212EF9),
   .weight23_1_pe5(24'h2532D7),
   .weight24_1_pe5(24'hFEBF15),
   .weight25_1_pe5(24'hD8F1EB),
   .weight26_1_pe5(24'h477FF1),
   .weight27_1_pe5(24'h304A19),
   .weight28_1_pe5(24'h3F0511),
   .weight29_1_pe5(24'hF6320C),
   .weight30_1_pe5(24'h2CE62A),
   .weight31_1_pe5(24'h26005E),
   .weight32_1_pe5(24'hD9D1BE),
   .weight33_1_pe5(24'h443A44),
   .weight34_1_pe5(24'hB47CEF),
   .weight35_1_pe5(24'h167F52),
   .weight36_1_pe5(24'h183F97),
   .weight01_2_pe5(24'hF50C5F),
   .weight02_2_pe5(24'h18F73E),
   .weight03_2_pe5(24'h0AE62C),
   .weight04_2_pe5(24'hD6B87C),
   .weight05_2_pe5(24'hFF7932),
   .weight06_2_pe5(24'h24C5D5),
   .weight07_2_pe5(24'h2BB0CA),
   .weight08_2_pe5(24'h6F7FF7),
   .weight09_2_pe5(24'h132C24),
   .weight10_2_pe5(24'h731EC9),
   .weight11_2_pe5(24'h036D06),
   .weight12_2_pe5(24'hFD120C),
   .weight13_2_pe5(24'hE00B35),
   .weight14_2_pe5(24'hCC7F37),
   .weight15_2_pe5(24'h3B204E),
   .weight16_2_pe5(24'h7F97B6),
   .weight17_2_pe5(24'h465F4B),
   .weight18_2_pe5(24'hE8F3DB),
   .weight19_2_pe5(24'h6E4D68),
   .weight20_2_pe5(24'hEE3B05),
   .weight21_2_pe5(24'h7E4FED),
   .weight22_2_pe5(24'hC2A98F),
   .weight23_2_pe5(24'hE211B6),
   .weight24_2_pe5(24'h00BAFB),
   .weight25_2_pe5(24'h877F67),
   .weight26_2_pe5(24'hA17F80),
   .weight27_2_pe5(24'hDBF200),
   .weight28_2_pe5(24'h090EF5),
   .weight29_2_pe5(24'hFE7F80),
   .weight30_2_pe5(24'hAF0085),
   .weight31_2_pe5(24'hC6B996),
   .weight32_2_pe5(24'hCA7FC3),
   .weight33_2_pe5(24'hBFEBF1),
   .weight34_2_pe5(24'hB93F14),
   .weight35_2_pe5(24'h2A2FC9),
   .weight36_2_pe5(24'h200B41)
)core_layer2(
   .i_clk(i_clk),
   .i_rstn(i_rstn),
   .s_axis_tready(m_axis_tready_core[0]),
   .s_axis_tvalid(m_axis_tvalid_core[0]),
   .s_axis_tdata(m_axis_tdata_core[0]),
   .m_axis_tdata(m_axis_tdata_core[1]),
   .m_axis_tvalid(m_axis_tvalid_core[1]),
   .m_axis_tready(m_axis_tready_core[1]),
   .EOL(),
   .EOF()
);

Axi4ConvCore#(
   .REQUANT(55),
   .weight01_1_pe0(24'h5B377F),
   .weight02_1_pe0(24'h074290),
   .weight03_1_pe0(24'h0ECCB4),
   .weight04_1_pe0(24'hF7F3FE),
   .weight05_1_pe0(24'hFDF7F7),
   .weight06_1_pe0(24'hFE0DF9),
   .weight07_1_pe0(24'hE224B9),
   .weight08_1_pe0(24'h807FEB),
   .weight09_1_pe0(24'h0F13E2),
   .weight10_1_pe0(24'h3FA234),
   .weight11_1_pe0(24'h376D23),
   .weight12_1_pe0(24'h854808),
   .weight13_1_pe0(24'h113CFC),
   .weight14_1_pe0(24'hE47F5D),
   .weight15_1_pe0(24'h2DE71D),
   .weight16_1_pe0(24'h1F622B),
   .weight17_1_pe0(24'h157F31),
   .weight18_1_pe0(24'h1F4615),
   .weight19_1_pe0(24'hC99B20),
   .weight20_1_pe0(24'h0C6CAD),
   .weight21_1_pe0(24'hBF0637),
   .weight22_1_pe0(24'hEDC92D),
   .weight23_1_pe0(24'h487FED),
   .weight24_1_pe0(24'hC548E0),
   .weight25_1_pe0(24'hF2AB38),
   .weight26_1_pe0(24'hA17FD5),
   .weight27_1_pe0(24'hE027F5),
   .weight28_1_pe0(24'h4F67D1),
   .weight29_1_pe0(24'hB2F183),
   .weight30_1_pe0(24'h1BA9DE),
   .weight31_1_pe0(24'hB327FD),
   .weight32_1_pe0(24'h417F1C),
   .weight33_1_pe0(24'h14F847),
   .weight34_1_pe0(24'hDF8C7D),
   .weight35_1_pe0(24'h434902),
   .weight36_1_pe0(24'hC705B5),
   .weight01_2_pe0(24'h1A8098),
   .weight02_2_pe0(24'hD87992),
   .weight03_2_pe0(24'h12D711),
   .weight04_2_pe0(24'hECFCF1),
   .weight05_2_pe0(24'hEC0EF4),
   .weight06_2_pe0(24'h09F20C),
   .weight07_2_pe0(24'h1A09DF),
   .weight08_2_pe0(24'h177F4C),
   .weight09_2_pe0(24'h04D6D6),
   .weight10_2_pe0(24'h7FFEFB),
   .weight11_2_pe0(24'hD97F38),
   .weight12_2_pe0(24'hBB5773),
   .weight13_2_pe0(24'h7A7F4D),
   .weight14_2_pe0(24'h05067E),
   .weight15_2_pe0(24'hE04D08),
   .weight16_2_pe0(24'hFAD081),
   .weight17_2_pe0(24'h7FE525),
   .weight18_2_pe0(24'hF20234),
   .weight19_2_pe0(24'h097F58),
   .weight20_2_pe0(24'hB97F4E),
   .weight21_2_pe0(24'hF8D7EE),
   .weight22_2_pe0(24'hFC000C),
   .weight23_2_pe0(24'hEEA6DF),
   .weight24_2_pe0(24'h11C334),
   .weight25_2_pe0(24'h195411),
   .weight26_2_pe0(24'h68B8E7),
   .weight27_2_pe0(24'h6007CD),
   .weight28_2_pe0(24'hEA46C0),
   .weight29_2_pe0(24'h827FE4),
   .weight30_2_pe0(24'hD338D8),
   .weight31_2_pe0(24'hEADE21),
   .weight32_2_pe0(24'hEB8014),
   .weight33_2_pe0(24'hF9DDEE),
   .weight34_2_pe0(24'h10E0FE),
   .weight35_2_pe0(24'hFE80C4),
   .weight36_2_pe0(24'hF2251A),
   .weight01_1_pe1(24'hF0280D),
   .weight02_1_pe1(24'hD840F9),
   .weight03_1_pe1(24'h18E3CE),
   .weight04_1_pe1(24'hFC0A03),
   .weight05_1_pe1(24'hFD00EE),
   .weight06_1_pe1(24'hEE00F3),
   .weight07_1_pe1(24'hFD41E3),
   .weight08_1_pe1(24'h155679),
   .weight09_1_pe1(24'h4FFAEB),
   .weight10_1_pe1(24'hF32628),
   .weight11_1_pe1(24'h7F7F0E),
   .weight12_1_pe1(24'h6F1703),
   .weight13_1_pe1(24'h2C38EE),
   .weight14_1_pe1(24'h9F7FF5),
   .weight15_1_pe1(24'h9C3E55),
   .weight16_1_pe1(24'hE9812F),
   .weight17_1_pe1(24'h172BE3),
   .weight18_1_pe1(24'h4D783E),
   .weight19_1_pe1(24'h0656F7),
   .weight20_1_pe1(24'h814B71),
   .weight21_1_pe1(24'h1A02D2),
   .weight22_1_pe1(24'h81D817),
   .weight23_1_pe1(24'h986ABE),
   .weight24_1_pe1(24'h7302F1),
   .weight25_1_pe1(24'hFF338C),
   .weight26_1_pe1(24'h8C7FA7),
   .weight27_1_pe1(24'h6B9CE6),
   .weight28_1_pe1(24'h137F00),
   .weight29_1_pe1(24'h953F5E),
   .weight30_1_pe1(24'hBCB910),
   .weight31_1_pe1(24'h35D5F3),
   .weight32_1_pe1(24'hD07F0B),
   .weight33_1_pe1(24'hCC81EB),
   .weight34_1_pe1(24'h9513E2),
   .weight35_1_pe1(24'h800C4D),
   .weight36_1_pe1(24'hE2060D),
   .weight01_2_pe1(24'h4580F1),
   .weight02_2_pe1(24'h016F7F),
   .weight03_2_pe1(24'h141F40),
   .weight04_2_pe1(24'h04F4F7),
   .weight05_2_pe1(24'h0B09F4),
   .weight06_2_pe1(24'hF814F6),
   .weight07_2_pe1(24'hEED02D),
   .weight08_2_pe1(24'h160EC7),
   .weight09_2_pe1(24'hD88019),
   .weight10_2_pe1(24'hD931FC),
   .weight11_2_pe1(24'h7F80CD),
   .weight12_2_pe1(24'hCAF380),
   .weight13_2_pe1(24'hE7FFF9),
   .weight14_2_pe1(24'hDB7F0B),
   .weight15_2_pe1(24'hDB38D5),
   .weight16_2_pe1(24'hF434F2),
   .weight17_2_pe1(24'h157F0B),
   .weight18_2_pe1(24'h192FEE),
   .weight19_2_pe1(24'hD201DA),
   .weight20_2_pe1(24'h183DD4),
   .weight21_2_pe1(24'h1422ED),
   .weight22_2_pe1(24'h06FB07),
   .weight23_2_pe1(24'hE77FD1),
   .weight24_2_pe1(24'hFD7216),
   .weight25_2_pe1(24'h0831D6),
   .weight26_2_pe1(24'h087F2E),
   .weight27_2_pe1(24'h0755FA),
   .weight28_2_pe1(24'h23EB29),
   .weight29_2_pe1(24'h472F30),
   .weight30_2_pe1(24'h0AE41A),
   .weight31_2_pe1(24'h04F943),
   .weight32_2_pe1(24'hD67FE5),
   .weight33_2_pe1(24'hCE5BF5),
   .weight34_2_pe1(24'h0016E5),
   .weight35_2_pe1(24'h287929),
   .weight36_2_pe1(24'h3F0B1D),
   .weight01_1_pe2(24'hD680BD),
   .weight02_1_pe2(24'h296780),
   .weight03_1_pe2(24'hF1D8D5),
   .weight04_1_pe2(24'h0B0AFB),
   .weight05_1_pe2(24'hFA06F3),
   .weight06_1_pe2(24'h04F20B),
   .weight07_1_pe2(24'h0FF02D),
   .weight08_1_pe2(24'h22041B),
   .weight09_1_pe2(24'h201D02),
   .weight10_1_pe2(24'h395AE6),
   .weight11_1_pe2(24'h2C7FB7),
   .weight12_1_pe2(24'h45923B),
   .weight13_1_pe2(24'h1709FC),
   .weight14_1_pe2(24'h4C7FCF),
   .weight15_1_pe2(24'hD70272),
   .weight16_1_pe2(24'h5C4813),
   .weight17_1_pe2(24'hF17F1F),
   .weight18_1_pe2(24'h01214E),
   .weight19_1_pe2(24'h153617),
   .weight20_1_pe2(24'h227EFE),
   .weight21_1_pe2(24'h1BD9E3),
   .weight22_1_pe2(24'hF718E5),
   .weight23_1_pe2(24'h507FA7),
   .weight24_1_pe2(24'h35AD1A),
   .weight25_1_pe2(24'h0F37F8),
   .weight26_1_pe2(24'hB07FC7),
   .weight27_1_pe2(24'hFADE11),
   .weight28_1_pe2(24'h99094D),
   .weight29_1_pe2(24'hC94860),
   .weight30_1_pe2(24'hFBF4F2),
   .weight31_1_pe2(24'h01E1B8),
   .weight32_1_pe2(24'h6F7FEA),
   .weight33_1_pe2(24'h1F07EC),
   .weight34_1_pe2(24'hDE21E5),
   .weight35_1_pe2(24'hA67FAF),
   .weight36_1_pe2(24'hECE4F4),
   .weight01_2_pe2(24'hFB07DE),
   .weight02_2_pe2(24'h22C147),
   .weight03_2_pe2(24'hAF33EE),
   .weight04_2_pe2(24'hFCF8F2),
   .weight05_2_pe2(24'h140A11),
   .weight06_2_pe2(24'hFF0106),
   .weight07_2_pe2(24'h0210D4),
   .weight08_2_pe2(24'hEC37FD),
   .weight09_2_pe2(24'hBA0720),
   .weight10_2_pe2(24'hB8DE1B),
   .weight11_2_pe2(24'h9202CC),
   .weight12_2_pe2(24'h957F00),
   .weight13_2_pe2(24'hE3DE06),
   .weight14_2_pe2(24'h307FE5),
   .weight15_2_pe2(24'hE8E201),
   .weight16_2_pe2(24'h18361D),
   .weight17_2_pe2(24'h377EF8),
   .weight18_2_pe2(24'h00BE02),
   .weight19_2_pe2(24'hC7011E),
   .weight20_2_pe2(24'hD17FAC),
   .weight21_2_pe2(24'hEA1AF1),
   .weight22_2_pe2(24'h5230FE),
   .weight23_2_pe2(24'h407F43),
   .weight24_2_pe2(24'hE408CE),
   .weight25_2_pe2(24'h213103),
   .weight26_2_pe2(24'h2D7F26),
   .weight27_2_pe2(24'h1A32FB),
   .weight28_2_pe2(24'hE68611),
   .weight29_2_pe2(24'h10260E),
   .weight30_2_pe2(24'h0119F5),
   .weight31_2_pe2(24'h2459C4),
   .weight32_2_pe2(24'h757F35),
   .weight33_2_pe2(24'h041EFA),
   .weight34_2_pe2(24'h15CCFF),
   .weight35_2_pe2(24'h2956F3),
   .weight36_2_pe2(24'hF600DF),
   .weight01_1_pe3(24'hC165F3),
   .weight02_1_pe3(24'h137F05),
   .weight03_1_pe3(24'h04D6F6),
   .weight04_1_pe3(24'h01EE10),
   .weight05_1_pe3(24'hFC04FD),
   .weight06_1_pe3(24'hF6F808),
   .weight07_1_pe3(24'h3E62BA),
   .weight08_1_pe3(24'h05429A),
   .weight09_1_pe3(24'hC5DC9A),
   .weight10_1_pe3(24'hDAE756),
   .weight11_1_pe3(24'h7F801C),
   .weight12_1_pe3(24'h458023),
   .weight13_1_pe3(24'hDF5375),
   .weight14_1_pe3(24'h46F855),
   .weight15_1_pe3(24'hCD075C),
   .weight16_1_pe3(24'h9E9D8A),
   .weight17_1_pe3(24'h28DC81),
   .weight18_1_pe3(24'h427F3C),
   .weight19_1_pe3(24'hA5EF34),
   .weight20_1_pe3(24'h69EB7F),
   .weight21_1_pe3(24'h3EF7F4),
   .weight22_1_pe3(24'h1F7F78),
   .weight23_1_pe3(24'h03AD81),
   .weight24_1_pe3(24'hF5C443),
   .weight25_1_pe3(24'h43DAB8),
   .weight26_1_pe3(24'h7F5F06),
   .weight27_1_pe3(24'h7F5893),
   .weight28_1_pe3(24'hE86295),
   .weight29_1_pe3(24'h9787B5),
   .weight30_1_pe3(24'hADE3E7),
   .weight31_1_pe3(24'h22511B),
   .weight32_1_pe3(24'hC7236C),
   .weight33_1_pe3(24'h86FCFB),
   .weight34_1_pe3(24'hE48EFA),
   .weight35_1_pe3(24'h07817F),
   .weight36_1_pe3(24'h38F27F),
   .weight01_2_pe3(24'hFE0010),
   .weight02_2_pe3(24'h09EEFA),
   .weight03_2_pe3(24'h03EDF8),
   .weight04_2_pe3(24'h05F3FE),
   .weight05_2_pe3(24'hFCF2FF),
   .weight06_2_pe3(24'h090CFF),
   .weight07_2_pe3(24'hF6F0FF),
   .weight08_2_pe3(24'hF4EF00),
   .weight09_2_pe3(24'hEDEB08),
   .weight10_2_pe3(24'hF10B0F),
   .weight11_2_pe3(24'hFFE9F3),
   .weight12_2_pe3(24'hF7EDF4),
   .weight13_2_pe3(24'h07F105),
   .weight14_2_pe3(24'hF9F2FC),
   .weight15_2_pe3(24'h01ED08),
   .weight16_2_pe3(24'h06F00C),
   .weight17_2_pe3(24'hFCF7F0),
   .weight18_2_pe3(24'hFD00F5),
   .weight19_2_pe3(24'hEF09F5),
   .weight20_2_pe3(24'h0C07F3),
   .weight21_2_pe3(24'hEEEEEE),
   .weight22_2_pe3(24'hFB05ED),
   .weight23_2_pe3(24'hF205FF),
   .weight24_2_pe3(24'h0DEE0F),
   .weight25_2_pe3(24'hECFEF4),
   .weight26_2_pe3(24'hFF0609),
   .weight27_2_pe3(24'h03F5ED),
   .weight28_2_pe3(24'h11F7FD),
   .weight29_2_pe3(24'h01FD0B),
   .weight30_2_pe3(24'hF6060E),
   .weight31_2_pe3(24'hF2F2FF),
   .weight32_2_pe3(24'hF200F7),
   .weight33_2_pe3(24'h09FF09),
   .weight34_2_pe3(24'h0A03FD),
   .weight35_2_pe3(24'h04EEF7),
   .weight36_2_pe3(24'hF9E7EE),
   .weight01_1_pe4(24'hEB34F6),
   .weight02_1_pe4(24'h1076AA),
   .weight03_1_pe4(24'hBDE523),
   .weight04_1_pe4(24'hF90E08),
   .weight05_1_pe4(24'h08040E),
   .weight06_1_pe4(24'hF5F712),
   .weight07_1_pe4(24'h0411F5),
   .weight08_1_pe4(24'h087FA4),
   .weight09_1_pe4(24'hC1FE19),
   .weight10_1_pe4(24'h6E7926),
   .weight11_1_pe4(24'h176064),
   .weight12_1_pe4(24'hE27B3D),
   .weight13_1_pe4(24'hDEB84E),
   .weight14_1_pe4(24'h7F8118),
   .weight15_1_pe4(24'h53436F),
   .weight16_1_pe4(24'h7F77D5),
   .weight17_1_pe4(24'h7F7F2F),
   .weight18_1_pe4(24'hD773E2),
   .weight19_1_pe4(24'hC31127),
   .weight20_1_pe4(24'h2D59DF),
   .weight21_1_pe4(24'h80A833),
   .weight22_1_pe4(24'hC38E15),
   .weight23_1_pe4(24'hF180E8),
   .weight24_1_pe4(24'h868223),
   .weight25_1_pe4(24'h280FBB),
   .weight26_1_pe4(24'h7F815C),
   .weight27_1_pe4(24'h1608E4),
   .weight28_1_pe4(24'hD6DEE7),
   .weight29_1_pe4(24'hAD21CD),
   .weight30_1_pe4(24'h2649C8),
   .weight31_1_pe4(24'h01444A),
   .weight32_1_pe4(24'h5081E2),
   .weight33_1_pe4(24'h0443DE),
   .weight34_1_pe4(24'hF2CA26),
   .weight35_1_pe4(24'h7F82C7),
   .weight36_1_pe4(24'hFF1CD3),
   .weight01_2_pe4(24'hAD32EF),
   .weight02_2_pe4(24'h11B7EC),
   .weight03_2_pe4(24'hFEA90A),
   .weight04_2_pe4(24'hFD1705),
   .weight05_2_pe4(24'h05FBF8),
   .weight06_2_pe4(24'hF0FCF7),
   .weight07_2_pe4(24'h415EB2),
   .weight08_2_pe4(24'h208068),
   .weight09_2_pe4(24'hF310D3),
   .weight10_2_pe4(24'hA6F958),
   .weight11_2_pe4(24'h7F6E5F),
   .weight12_2_pe4(24'h6C807F),
   .weight13_2_pe4(24'hD81AF6),
   .weight14_2_pe4(24'hD77F5F),
   .weight15_2_pe4(24'h117A20),
   .weight16_2_pe4(24'h086C02),
   .weight17_2_pe4(24'hBD7F5F),
   .weight18_2_pe4(24'hFC7D3C),
   .weight19_2_pe4(24'h274B54),
   .weight20_2_pe4(24'h602F7F),
   .weight21_2_pe4(24'h08C8FA),
   .weight22_2_pe4(24'hAACAF5),
   .weight23_2_pe4(24'hCF7FE1),
   .weight24_2_pe4(24'h0DB81B),
   .weight25_2_pe4(24'h38EDCE),
   .weight26_2_pe4(24'h267F24),
   .weight27_2_pe4(24'h10E230),
   .weight28_2_pe4(24'h16E4D9),
   .weight29_2_pe4(24'h7FE18C),
   .weight30_2_pe4(24'h0A0CCC),
   .weight31_2_pe4(24'h37BD18),
   .weight32_2_pe4(24'hF47F38),
   .weight33_2_pe4(24'hEDCE1A),
   .weight34_2_pe4(24'hA41411),
   .weight35_2_pe4(24'h947FDC),
   .weight36_2_pe4(24'h11C800),
   .weight01_1_pe5(24'h0C01F9),
   .weight02_1_pe5(24'h080CF7),
   .weight03_1_pe5(24'hF805F6),
   .weight04_1_pe5(24'h04F902),
   .weight05_1_pe5(24'hF6100C),
   .weight06_1_pe5(24'h0E0203),
   .weight07_1_pe5(24'hF5EDF4),
   .weight08_1_pe5(24'hFA02F8),
   .weight09_1_pe5(24'h00F209),
   .weight10_1_pe5(24'hFEF8EE),
   .weight11_1_pe5(24'h09E6ED),
   .weight12_1_pe5(24'hF8EB0B),
   .weight13_1_pe5(24'hF0F301),
   .weight14_1_pe5(24'hFF0C0E),
   .weight15_1_pe5(24'hFAEDFB),
   .weight16_1_pe5(24'h04F008),
   .weight17_1_pe5(24'hF0F20D),
   .weight18_1_pe5(24'h0502F2),
   .weight19_1_pe5(24'hF000F3),
   .weight20_1_pe5(24'hFCEBF2),
   .weight21_1_pe5(24'h0EE3FB),
   .weight22_1_pe5(24'hECFEFC),
   .weight23_1_pe5(24'h04E9F7),
   .weight24_1_pe5(24'h070707),
   .weight25_1_pe5(24'hFFF5FC),
   .weight26_1_pe5(24'h08F6EA),
   .weight27_1_pe5(24'hEDF80B),
   .weight28_1_pe5(24'h0D02F2),
   .weight29_1_pe5(24'h04E8EA),
   .weight30_1_pe5(24'hEEFDFD),
   .weight31_1_pe5(24'hEC0A0A),
   .weight32_1_pe5(24'h00E9EB),
   .weight33_1_pe5(24'h00FDF6),
   .weight34_1_pe5(24'h08ECF8),
   .weight35_1_pe5(24'hF90C0F),
   .weight36_1_pe5(24'hF001FD),
   .weight01_2_pe5(24'h9F5FF3),
   .weight02_2_pe5(24'hE7802F),
   .weight03_2_pe5(24'h3D4325),
   .weight04_2_pe5(24'hF707F9),
   .weight05_2_pe5(24'hF0F210),
   .weight06_2_pe5(24'hF8F802),
   .weight07_2_pe5(24'h08C641),
   .weight08_2_pe5(24'h639BB4),
   .weight09_2_pe5(24'h1569FA),
   .weight10_2_pe5(24'h2600C9),
   .weight11_2_pe5(24'h819B43),
   .weight12_2_pe5(24'h7F27D9),
   .weight13_2_pe5(24'hE628F8),
   .weight14_2_pe5(24'h727F30),
   .weight15_2_pe5(24'hB9FFCD),
   .weight16_2_pe5(24'hD12C0F),
   .weight17_2_pe5(24'hE87FFE),
   .weight18_2_pe5(24'h06DDF5),
   .weight19_2_pe5(24'h4CF0FE),
   .weight20_2_pe5(24'h116519),
   .weight21_2_pe5(24'h341F24),
   .weight22_2_pe5(24'h151CC2),
   .weight23_2_pe5(24'hFC7F0B),
   .weight24_2_pe5(24'h6312F6),
   .weight25_2_pe5(24'hB4EEFC),
   .weight26_2_pe5(24'hF57F31),
   .weight27_2_pe5(24'h1701BC),
   .weight28_2_pe5(24'h1106ED),
   .weight29_2_pe5(24'hBF33EF),
   .weight30_2_pe5(24'hED5005),
   .weight31_2_pe5(24'h26262C),
   .weight32_2_pe5(24'hEE7F06),
   .weight33_2_pe5(24'hFF3014),
   .weight34_2_pe5(24'hE3E427),
   .weight35_2_pe5(24'hD97F16),
   .weight36_2_pe5(24'hF0F538)
)core_layer3(
   .i_clk(i_clk),
   .i_rstn(i_rstn),
   .s_axis_tready(m_axis_tready_core[1]),
   .s_axis_tvalid(m_axis_tvalid_core[1]),
   .s_axis_tdata(m_axis_tdata_core[1]),
   .m_axis_tdata(m_axis_tdata_core[2]),
   .m_axis_tvalid(m_axis_tvalid_core[2]),
   .m_axis_tready(m_axis_tready_core[2]),
   .EOL(),
   .EOF()
);

Axi4ConvCore#(
   .REQUANT(109),
   .weight01_1_pe0(24'h0CFB01),
   .weight02_1_pe0(24'h0C09EF),
   .weight03_1_pe0(24'h10EFEB),
   .weight04_1_pe0(24'hF102E8),
   .weight05_1_pe0(24'hEEFDF0),
   .weight06_1_pe0(24'hECF30F),
   .weight07_1_pe0(24'hE9E8E2),
   .weight08_1_pe0(24'hEC050F),
   .weight09_1_pe0(24'hFCED07),
   .weight10_1_pe0(24'hF5F4F8),
   .weight11_1_pe0(24'h0C150E),
   .weight12_1_pe0(24'hE5FD12),
   .weight13_1_pe0(24'hE4DCEA),
   .weight14_1_pe0(24'hF600F2),
   .weight15_1_pe0(24'h09ECE4),
   .weight16_1_pe0(24'h1D0C1A),
   .weight17_1_pe0(24'h110714),
   .weight18_1_pe0(24'hFAF9FB),
   .weight19_1_pe0(24'hF1FEF5),
   .weight20_1_pe0(24'hFAF7F9),
   .weight21_1_pe0(24'hE9E5DE),
   .weight22_1_pe0(24'hE4FF11),
   .weight23_1_pe0(24'h15DCDF),
   .weight24_1_pe0(24'h07F113),
   .weight25_1_pe0(24'hED05E0),
   .weight26_1_pe0(24'hE90AE6),
   .weight27_1_pe0(24'hE91105),
   .weight28_1_pe0(24'h0504EE),
   .weight29_1_pe0(24'h01EEED),
   .weight30_1_pe0(24'h0B04EE),
   .weight31_1_pe0(24'h160F00),
   .weight32_1_pe0(24'hF6F8E6),
   .weight33_1_pe0(24'h08060F),
   .weight34_1_pe0(24'hF3DB09),
   .weight35_1_pe0(24'hFF04F4),
   .weight36_1_pe0(24'hED03ED),
   .weight01_2_pe0(24'hEC9BED),
   .weight02_2_pe0(24'h097FBE),
   .weight03_2_pe0(24'hD9091E),
   .weight04_2_pe0(24'hF4A7F3),
   .weight05_2_pe0(24'hFE7C91),
   .weight06_2_pe0(24'h1FE312),
   .weight07_2_pe0(24'h0AE113),
   .weight08_2_pe0(24'h4E7F11),
   .weight09_2_pe0(24'h0805EA),
   .weight10_2_pe0(24'h1CF90F),
   .weight11_2_pe0(24'hE33F6A),
   .weight12_2_pe0(24'h090AFC),
   .weight13_2_pe0(24'h024105),
   .weight14_2_pe0(24'h09C322),
   .weight15_2_pe0(24'hF938D7),
   .weight16_2_pe0(24'hE904F5),
   .weight17_2_pe0(24'h15E9E2),
   .weight18_2_pe0(24'h1100FD),
   .weight19_2_pe0(24'hDC5213),
   .weight20_2_pe0(24'h2528FF),
   .weight21_2_pe0(24'hB5C108),
   .weight22_2_pe0(24'h384310),
   .weight23_2_pe0(24'hEF6FCB),
   .weight24_2_pe0(24'h10E011),
   .weight25_2_pe0(24'hE1B5CF),
   .weight26_2_pe0(24'h017F10),
   .weight27_2_pe0(24'h1E19F0),
   .weight28_2_pe0(24'h1EE5EB),
   .weight29_2_pe0(24'hE9EA06),
   .weight30_2_pe0(24'hF6FF08),
   .weight31_2_pe0(24'hC2BD24),
   .weight32_2_pe0(24'h7F6A19),
   .weight33_2_pe0(24'hDA1EEB),
   .weight34_2_pe0(24'hE2F506),
   .weight35_2_pe0(24'h07123B),
   .weight36_2_pe0(24'hD726F6),
   .weight01_1_pe1(24'h808080),
   .weight02_1_pe1(24'h517D25),
   .weight03_1_pe1(24'hE9CFED),
   .weight04_1_pe1(24'h808080),
   .weight05_1_pe1(24'hDE8046),
   .weight06_1_pe1(24'h03561F),
   .weight07_1_pe1(24'h808080),
   .weight08_1_pe1(24'h8072FB),
   .weight09_1_pe1(24'h5DCDAC),
   .weight10_1_pe1(24'h808080),
   .weight11_1_pe1(24'h6507F7),
   .weight12_1_pe1(24'hCC4F08),
   .weight13_1_pe1(24'h808080),
   .weight14_1_pe1(24'h167F0A),
   .weight15_1_pe1(24'hF6BDD9),
   .weight16_1_pe1(24'hEAE6E7),
   .weight17_1_pe1(24'h080101),
   .weight18_1_pe1(24'h01F901),
   .weight19_1_pe1(24'h808080),
   .weight20_1_pe1(24'hBE80FE),
   .weight21_1_pe1(24'h3B7FA6),
   .weight22_1_pe1(24'h808080),
   .weight23_1_pe1(24'h087D01),
   .weight24_1_pe1(24'h122DFC),
   .weight25_1_pe1(24'h808080),
   .weight26_1_pe1(24'hEF7FD4),
   .weight27_1_pe1(24'h1713F1),
   .weight28_1_pe1(24'h16F4F7),
   .weight29_1_pe1(24'h1A12DC),
   .weight30_1_pe1(24'hFAFF16),
   .weight31_1_pe1(24'h808080),
   .weight32_1_pe1(24'h912C52),
   .weight33_1_pe1(24'h0430FD),
   .weight34_1_pe1(24'h808080),
   .weight35_1_pe1(24'h117F43),
   .weight36_1_pe1(24'hC0ACFC),
   .weight01_2_pe1(24'hB3FC34),
   .weight02_2_pe1(24'h2D3449),
   .weight03_2_pe1(24'hF571E8),
   .weight04_2_pe1(24'h33805E),
   .weight05_2_pe1(24'hF3207F),
   .weight06_2_pe1(24'hF4CB02),
   .weight07_2_pe1(24'hA74ACE),
   .weight08_2_pe1(24'h2338E4),
   .weight09_2_pe1(24'h08860D),
   .weight10_2_pe1(24'h507FE6),
   .weight11_2_pe1(24'hE47FD4),
   .weight12_2_pe1(24'h0D2CD7),
   .weight13_2_pe1(24'hCC7ECC),
   .weight14_2_pe1(24'h568480),
   .weight15_2_pe1(24'h3BD533),
   .weight16_2_pe1(24'h0817FE),
   .weight17_2_pe1(24'h0C0A10),
   .weight18_2_pe1(24'hF4EAF6),
   .weight19_2_pe1(24'h245CB1),
   .weight20_2_pe1(24'h7F56DE),
   .weight21_2_pe1(24'h019FC6),
   .weight22_2_pe1(24'hE05DD8),
   .weight23_2_pe1(24'hC67FD4),
   .weight24_2_pe1(24'h20B6FE),
   .weight25_2_pe1(24'h682572),
   .weight26_2_pe1(24'h1C2676),
   .weight27_2_pe1(24'hE321D1),
   .weight28_2_pe1(24'h0419F5),
   .weight29_2_pe1(24'h06080E),
   .weight30_2_pe1(24'h130B0C),
   .weight31_2_pe1(24'h9740EB),
   .weight32_2_pe1(24'hC97FFE),
   .weight33_2_pe1(24'hCDFC49),
   .weight34_2_pe1(24'hE8F4A9),
   .weight35_2_pe1(24'hEE7FF6),
   .weight36_2_pe1(24'h23651D),
   .weight01_1_pe2(24'hD9BBEF),
   .weight02_1_pe2(24'h637F72),
   .weight03_1_pe2(24'h62AC86),
   .weight04_1_pe2(24'h1AF5D3),
   .weight05_1_pe2(24'h087F7F),
   .weight06_1_pe2(24'hA89A2C),
   .weight07_1_pe2(24'hAF823D),
   .weight08_1_pe2(24'h807F16),
   .weight09_1_pe2(24'hC57E3A),
   .weight10_1_pe2(24'hD6809E),
   .weight11_1_pe2(24'h8080B2),
   .weight12_1_pe2(24'h1080EE),
   .weight13_1_pe2(24'hE34859),
   .weight14_1_pe2(24'hCBBC94),
   .weight15_1_pe2(24'h0FFD62),
   .weight16_1_pe2(24'hFBF5E5),
   .weight17_1_pe2(24'h1EECEC),
   .weight18_1_pe2(24'h16F710),
   .weight19_1_pe2(24'h513127),
   .weight20_1_pe2(24'h4B8012),
   .weight21_1_pe2(24'h0380D4),
   .weight22_1_pe2(24'h307F22),
   .weight23_1_pe2(24'h907FE5),
   .weight24_1_pe2(24'hF6D4C8),
   .weight25_1_pe2(24'h1D99DD),
   .weight26_1_pe2(24'h387F7F),
   .weight27_1_pe2(24'h804D3F),
   .weight28_1_pe2(24'h0FECF1),
   .weight29_1_pe2(24'hEA011C),
   .weight30_1_pe2(24'hFEEE12),
   .weight31_1_pe2(24'h3F8416),
   .weight32_1_pe2(24'hD27F80),
   .weight33_1_pe2(24'hFE9838),
   .weight34_1_pe2(24'h063DA9),
   .weight35_1_pe2(24'h127F99),
   .weight36_1_pe2(24'h557F16),
   .weight01_2_pe2(24'h8031BA),
   .weight02_2_pe2(24'h807FA8),
   .weight03_2_pe2(24'h80B72E),
   .weight04_2_pe2(24'h8024D2),
   .weight05_2_pe2(24'h8079E6),
   .weight06_2_pe2(24'h80F65B),
   .weight07_2_pe2(24'h802D49),
   .weight08_2_pe2(24'h807FE2),
   .weight09_2_pe2(24'h800FFC),
   .weight10_2_pe2(24'h80E832),
   .weight11_2_pe2(24'h80267F),
   .weight12_2_pe2(24'h80DB39),
   .weight13_2_pe2(24'h808035),
   .weight14_2_pe2(24'h808016),
   .weight15_2_pe2(24'h8061B2),
   .weight16_2_pe2(24'hE80F1A),
   .weight17_2_pe2(24'hE4EC17),
   .weight18_2_pe2(24'h010B14),
   .weight19_2_pe2(24'h80B60F),
   .weight20_2_pe2(24'h807F21),
   .weight21_2_pe2(24'h808009),
   .weight22_2_pe2(24'h80F1BF),
   .weight23_2_pe2(24'h807FE1),
   .weight24_2_pe2(24'h803C00),
   .weight25_2_pe2(24'h8014DD),
   .weight26_2_pe2(24'h807F0E),
   .weight27_2_pe2(24'h8003EF),
   .weight28_2_pe2(24'h170715),
   .weight29_2_pe2(24'hE91B14),
   .weight30_2_pe2(24'h08100E),
   .weight31_2_pe2(24'h808022),
   .weight32_2_pe2(24'h80FA5D),
   .weight33_2_pe2(24'h807FD1),
   .weight34_2_pe2(24'h80A93E),
   .weight35_2_pe2(24'h803D06),
   .weight36_2_pe2(24'h80BDC3),
   .weight01_1_pe3(24'h7F6F43),
   .weight02_1_pe3(24'h501FF2),
   .weight03_1_pe3(24'h13AEE3),
   .weight04_1_pe3(24'hB2BB7F),
   .weight05_1_pe3(24'hC080A7),
   .weight06_1_pe3(24'hE0A780),
   .weight07_1_pe3(24'hFB12D6),
   .weight08_1_pe3(24'h817F7F),
   .weight09_1_pe3(24'hEE5761),
   .weight10_1_pe3(24'hDDD8E3),
   .weight11_1_pe3(24'h8080CB),
   .weight12_1_pe3(24'h0E4BAE),
   .weight13_1_pe3(24'h8082FC),
   .weight14_1_pe3(24'h558066),
   .weight15_1_pe3(24'h61A880),
   .weight16_1_pe3(24'hEF0EF8),
   .weight17_1_pe3(24'hFB0113),
   .weight18_1_pe3(24'h1DF81A),
   .weight19_1_pe3(24'h3EA1E4),
   .weight20_1_pe3(24'h7FEE62),
   .weight21_1_pe3(24'h1A7F7F),
   .weight22_1_pe3(24'h00B836),
   .weight23_1_pe3(24'h80F8E1),
   .weight24_1_pe3(24'hCE01DD),
   .weight25_1_pe3(24'h80C6A6),
   .weight26_1_pe3(24'h8666A4),
   .weight27_1_pe3(24'hA30706),
   .weight28_1_pe3(24'h0AF00C),
   .weight29_1_pe3(24'hF7F4F5),
   .weight30_1_pe3(24'hEC05F7),
   .weight31_1_pe3(24'h6E778D),
   .weight32_1_pe3(24'h637F1D),
   .weight33_1_pe3(24'h5B7C02),
   .weight34_1_pe3(24'hE2D228),
   .weight35_1_pe3(24'hFE79FB),
   .weight36_1_pe3(24'h2DBCAD),
   .weight01_2_pe3(24'h0E6F0F),
   .weight02_2_pe3(24'hCB7F36),
   .weight03_2_pe3(24'h679726),
   .weight04_2_pe3(24'hCB7FDE),
   .weight05_2_pe3(24'h270AA3),
   .weight06_2_pe3(24'h07F495),
   .weight07_2_pe3(24'h7FA145),
   .weight08_2_pe3(24'hC77FFE),
   .weight09_2_pe3(24'hFF7701),
   .weight10_2_pe3(24'hC20B38),
   .weight11_2_pe3(24'h65807F),
   .weight12_2_pe3(24'hF60A19),
   .weight13_2_pe3(24'hCA8032),
   .weight14_2_pe3(24'hAE7F5D),
   .weight15_2_pe3(24'hD231C1),
   .weight16_2_pe3(24'hF7E214),
   .weight17_2_pe3(24'h11F010),
   .weight18_2_pe3(24'h10EF0D),
   .weight19_2_pe3(24'hDDD9D7),
   .weight20_2_pe3(24'hB97F1D),
   .weight21_2_pe3(24'h2EDB71),
   .weight22_2_pe3(24'h99ECBD),
   .weight23_2_pe3(24'h7FAFFC),
   .weight24_2_pe3(24'hEE1ECB),
   .weight25_2_pe3(24'hFC7FEC),
   .weight26_2_pe3(24'h287FB7),
   .weight27_2_pe3(24'hDEECF6),
   .weight28_2_pe3(24'h01F4FA),
   .weight29_2_pe3(24'hEF19E9),
   .weight30_2_pe3(24'hFC1613),
   .weight31_2_pe3(24'h7FA0BA),
   .weight32_2_pe3(24'h7F81D0),
   .weight33_2_pe3(24'h0CD3EB),
   .weight34_2_pe3(24'h0A330D),
   .weight35_2_pe3(24'h5F5D41),
   .weight36_2_pe3(24'h9C024E),
   .weight01_1_pe4(24'h364AE3),
   .weight02_1_pe4(24'hC842D0),
   .weight03_1_pe4(24'hF9EAFC),
   .weight04_1_pe4(24'hF34AD6),
   .weight05_1_pe4(24'h1380C5),
   .weight06_1_pe4(24'hFB4724),
   .weight07_1_pe4(24'h5B07D3),
   .weight08_1_pe4(24'hA27F32),
   .weight09_1_pe4(24'hFD46D2),
   .weight10_1_pe4(24'hC9ACE0),
   .weight11_1_pe4(24'hFE80C2),
   .weight12_1_pe4(24'hE2EF14),
   .weight13_1_pe4(24'h3EC718),
   .weight14_1_pe4(24'hCD7F36),
   .weight15_1_pe4(24'hFAECE4),
   .weight16_1_pe4(24'h001617),
   .weight17_1_pe4(24'h05F607),
   .weight18_1_pe4(24'hFD12F6),
   .weight19_1_pe4(24'hD28E33),
   .weight20_1_pe4(24'hAFB626),
   .weight21_1_pe4(24'h017F0D),
   .weight22_1_pe4(24'hF9FB06),
   .weight23_1_pe4(24'hFF7F24),
   .weight24_1_pe4(24'hF42D13),
   .weight25_1_pe4(24'hC11BE8),
   .weight26_1_pe4(24'h167F13),
   .weight27_1_pe4(24'h0BD74A),
   .weight28_1_pe4(24'hF7E108),
   .weight29_1_pe4(24'h0DF4EF),
   .weight30_1_pe4(24'h14FEEA),
   .weight31_1_pe4(24'h4935FB),
   .weight32_1_pe4(24'hC65BF8),
   .weight33_1_pe4(24'h34B8CB),
   .weight34_1_pe4(24'hFE1A18),
   .weight35_1_pe4(24'hF77F41),
   .weight36_1_pe4(24'h1D80CB),
   .weight01_2_pe4(24'h727FEE),
   .weight02_2_pe4(24'hA78A5B),
   .weight03_2_pe4(24'hF78BA9),
   .weight04_2_pe4(24'hF04AF2),
   .weight05_2_pe4(24'hF880CA),
   .weight06_2_pe4(24'h14302C),
   .weight07_2_pe4(24'h3887A3),
   .weight08_2_pe4(24'h91C630),
   .weight09_2_pe4(24'h5E4DF8),
   .weight10_2_pe4(24'h3164EC),
   .weight11_2_pe4(24'h0E80EB),
   .weight12_2_pe4(24'hA69508),
   .weight13_2_pe4(24'hFD8041),
   .weight14_2_pe4(24'hD57F35),
   .weight15_2_pe4(24'hEA9DB3),
   .weight16_2_pe4(24'hEEF619),
   .weight17_2_pe4(24'h1303E7),
   .weight18_2_pe4(24'h0DFFF0),
   .weight19_2_pe4(24'hC4802B),
   .weight20_2_pe4(24'hBF80D3),
   .weight21_2_pe4(24'h367412),
   .weight22_2_pe4(24'h4A7A72),
   .weight23_2_pe4(24'hF969E1),
   .weight24_2_pe4(24'hE73D1A),
   .weight25_2_pe4(24'hCE8B14),
   .weight26_2_pe4(24'h235584),
   .weight27_2_pe4(24'h05C86F),
   .weight28_2_pe4(24'h14F70F),
   .weight29_2_pe4(24'h11E4E8),
   .weight30_2_pe4(24'hF90B0E),
   .weight31_2_pe4(24'h61ADB5),
   .weight32_2_pe4(24'h821FE0),
   .weight33_2_pe4(24'h6BE545),
   .weight34_2_pe4(24'hD9C02F),
   .weight35_2_pe4(24'h166613),
   .weight36_2_pe4(24'h928581),
   .weight01_1_pe5(24'hC5FE26),
   .weight02_1_pe5(24'hC4943B),
   .weight03_1_pe5(24'h2F7F2E),
   .weight04_1_pe5(24'h094E50),
   .weight05_1_pe5(24'h7F7F31),
   .weight06_1_pe5(24'h05500A),
   .weight07_1_pe5(24'hFE09F8),
   .weight08_1_pe5(24'h7F80AF),
   .weight09_1_pe5(24'h358AEB),
   .weight10_1_pe5(24'h3D7A1B),
   .weight11_1_pe5(24'h7479DD),
   .weight12_1_pe5(24'hD40DDE),
   .weight13_1_pe5(24'h0BF3E1),
   .weight14_1_pe5(24'h0652C8),
   .weight15_1_pe5(24'hCFEFFC),
   .weight16_1_pe5(24'h180103),
   .weight17_1_pe5(24'hFA18F1),
   .weight18_1_pe5(24'h041802),
   .weight19_1_pe5(24'h0C19BA),
   .weight20_1_pe5(24'h0A7F03),
   .weight21_1_pe5(24'hF52428),
   .weight22_1_pe5(24'hDD9ADE),
   .weight23_1_pe5(24'h1CFF37),
   .weight24_1_pe5(24'h22EC2D),
   .weight25_1_pe5(24'h344561),
   .weight26_1_pe5(24'h4CA1CC),
   .weight27_1_pe5(24'h08F9B2),
   .weight28_1_pe5(24'h0119EA),
   .weight29_1_pe5(24'hE308FB),
   .weight30_1_pe5(24'h1907FB),
   .weight31_1_pe5(24'h04C8D3),
   .weight32_1_pe5(24'h80AD18),
   .weight33_1_pe5(24'hBCE1F9),
   .weight34_1_pe5(24'h0F18B3),
   .weight35_1_pe5(24'h16A9C8),
   .weight36_1_pe5(24'hD3EB16),
   .weight01_2_pe5(24'hDE001B),
   .weight02_2_pe5(24'h1F2F80),
   .weight03_2_pe5(24'hD55D80),
   .weight04_2_pe5(24'h3ACF80),
   .weight05_2_pe5(24'h0634F6),
   .weight06_2_pe5(24'h022F80),
   .weight07_2_pe5(24'hB67F80),
   .weight08_2_pe5(24'h8869A5),
   .weight09_2_pe5(24'h3F8080),
   .weight10_2_pe5(24'hFDEB80),
   .weight11_2_pe5(24'hCA7F80),
   .weight12_2_pe5(24'hF62080),
   .weight13_2_pe5(24'hFD32C5),
   .weight14_2_pe5(24'h01E480),
   .weight15_2_pe5(24'h17A580),
   .weight16_2_pe5(24'hEDEAED),
   .weight17_2_pe5(24'h0A05EC),
   .weight18_2_pe5(24'hE3F0F1),
   .weight19_2_pe5(24'h26CC80),
   .weight20_2_pe5(24'h628080),
   .weight21_2_pe5(24'h17A780),
   .weight22_2_pe5(24'h0BCFD5),
   .weight23_2_pe5(24'h0B7F80),
   .weight24_2_pe5(24'hFF1880),
   .weight25_2_pe5(24'h3CBA8E),
   .weight26_2_pe5(24'h655280),
   .weight27_2_pe5(24'h052E80),
   .weight28_2_pe5(24'hF60AFC),
   .weight29_2_pe5(24'hE310E8),
   .weight30_2_pe5(24'hFEF0E8),
   .weight31_2_pe5(24'hC95B80),
   .weight32_2_pe5(24'hDB7F2F),
   .weight33_2_pe5(24'hDDE780),
   .weight34_2_pe5(24'h160580),
   .weight35_2_pe5(24'hBD7F1C),
   .weight36_2_pe5(24'h02ED80)
)core_layer4(
   .i_clk(i_clk),
   .i_rstn(i_rstn),
   .s_axis_tready(m_axis_tready_core[2]),
   .s_axis_tvalid(m_axis_tvalid_core[2]),
   .s_axis_tdata(m_axis_tdata_core[2]),
   .m_axis_tdata(m_axis_tdata),
   .m_axis_tvalid(m_axis_tvalid),
   .m_axis_tready(m_axis_tready),
   .EOL(),
   .EOF()
);
   
endmodule